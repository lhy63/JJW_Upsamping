`timescale 1ns/1ps

module SuperResolutionCore (
  input               ddrDataIn_valid,
  output              ddrDataIn_ready,
  input      [31:0]   ddrDataIn_payload,
  input               ipConfig_aw_valid,
  output              ipConfig_aw_ready,
  input      [31:0]   ipConfig_aw_payload_addr,
  input      [2:0]    ipConfig_aw_payload_prot,
  input               ipConfig_w_valid,
  output              ipConfig_w_ready,
  input      [31:0]   ipConfig_w_payload_data,
  input      [3:0]    ipConfig_w_payload_strb,
  output              ipConfig_b_valid,
  input               ipConfig_b_ready,
  output     [1:0]    ipConfig_b_payload_resp,
  input               ipConfig_ar_valid,
  output              ipConfig_ar_ready,
  input      [31:0]   ipConfig_ar_payload_addr,
  input      [2:0]    ipConfig_ar_payload_prot,
  output              ipConfig_r_valid,
  input               ipConfig_r_ready,
  output     [31:0]   ipConfig_r_payload_data,
  output     [1:0]    ipConfig_r_payload_resp,
  output              inpDataOut_valid,
  input               inpDataOut_ready,
  output     [31:0]   inpDataOut_payload_pixel,
  output              inpDataOut_payload_frameStart,
  output              inpDataOut_payload_rowEnd,
  input               clk,
  input               resetn
);

  wire                ddrDataWrapper_1_ddrIn_ready;
  wire                ddrDataWrapper_1_pixelsOut_valid;
  wire       [31:0]   ddrDataWrapper_1_pixelsOut_payload_pixel;
  wire                ddrDataWrapper_1_pixelsOut_payload_frameStart;
  wire                ddrDataWrapper_1_pixelsOut_payload_rowEnd;
  wire                channelDispatcher_allPixelChannelIn_ready;
  wire                channelDispatcher_bPixelChannelOut_valid;
  wire       [7:0]    channelDispatcher_bPixelChannelOut_payload_pixel;
  wire                channelDispatcher_bPixelChannelOut_payload_frameStart;
  wire                channelDispatcher_bPixelChannelOut_payload_rowEnd;
  wire                channelDispatcher_gPixelChannelOut_valid;
  wire       [7:0]    channelDispatcher_gPixelChannelOut_payload_pixel;
  wire                channelDispatcher_gPixelChannelOut_payload_frameStart;
  wire                channelDispatcher_gPixelChannelOut_payload_rowEnd;
  wire                channelDispatcher_rPixelChannelOut_valid;
  wire       [7:0]    channelDispatcher_rPixelChannelOut_payload_pixel;
  wire                channelDispatcher_rPixelChannelOut_payload_frameStart;
  wire                channelDispatcher_rPixelChannelOut_payload_rowEnd;
  wire                bChannelPart1Core_pixelsIn_ready;
  wire                bChannelPart1Core_pixelsOut_valid;
  wire       [7:0]    bChannelPart1Core_pixelsOut_payload_pixel;
  wire                bChannelPart1Core_pixelsOut_payload_frameStart;
  wire                bChannelPart1Core_pixelsOut_payload_rowEnd;
  wire                bChannelPart1Core_startOut;
  wire                bChannelPart1Core_inpDoneOut;
  wire                bChannelPart2Core_pixelsIn_ready;
  wire                bChannelPart2Core_pixelsOut_valid;
  wire       [7:0]    bChannelPart2Core_pixelsOut_payload_pixel;
  wire                bChannelPart2Core_pixelsOut_payload_frameStart;
  wire                bChannelPart2Core_pixelsOut_payload_rowEnd;
  wire                bChannelPart2Core_pixelsOut_payload_inpValid;
  wire                bChannelPart2Core_startOut;
  wire                bChannelPart2Core_inpTwoDoneOut;
  wire                bChannelPart3Core_pixelsIn_ready;
  wire                bChannelPart3Core_pixelsOut_valid;
  wire       [7:0]    bChannelPart3Core_pixelsOut_payload_pixel;
  wire                bChannelPart3Core_pixelsOut_payload_frameStart;
  wire                bChannelPart3Core_pixelsOut_payload_rowEnd;
  wire                bChannelPart3Core_inpThreeDoneOut;
  wire                gChannelPart1Core_pixelsIn_ready;
  wire                gChannelPart1Core_pixelsOut_valid;
  wire       [7:0]    gChannelPart1Core_pixelsOut_payload_pixel;
  wire                gChannelPart1Core_pixelsOut_payload_frameStart;
  wire                gChannelPart1Core_pixelsOut_payload_rowEnd;
  wire                gChannelPart1Core_startOut;
  wire                gChannelPart1Core_inpDoneOut;
  wire                gChannelPart2Core_pixelsIn_ready;
  wire                gChannelPart2Core_pixelsOut_valid;
  wire       [7:0]    gChannelPart2Core_pixelsOut_payload_pixel;
  wire                gChannelPart2Core_pixelsOut_payload_frameStart;
  wire                gChannelPart2Core_pixelsOut_payload_rowEnd;
  wire                gChannelPart2Core_pixelsOut_payload_inpValid;
  wire                gChannelPart2Core_startOut;
  wire                gChannelPart2Core_inpTwoDoneOut;
  wire                gChannelPart3Core_pixelsIn_ready;
  wire                gChannelPart3Core_pixelsOut_valid;
  wire       [7:0]    gChannelPart3Core_pixelsOut_payload_pixel;
  wire                gChannelPart3Core_pixelsOut_payload_frameStart;
  wire                gChannelPart3Core_pixelsOut_payload_rowEnd;
  wire                gChannelPart3Core_inpThreeDoneOut;
  wire                rChannelPart1Core_pixelsIn_ready;
  wire                rChannelPart1Core_pixelsOut_valid;
  wire       [7:0]    rChannelPart1Core_pixelsOut_payload_pixel;
  wire                rChannelPart1Core_pixelsOut_payload_frameStart;
  wire                rChannelPart1Core_pixelsOut_payload_rowEnd;
  wire                rChannelPart1Core_startOut;
  wire                rChannelPart1Core_inpDoneOut;
  wire                rChannelPart2Core_pixelsIn_ready;
  wire                rChannelPart2Core_pixelsOut_valid;
  wire       [7:0]    rChannelPart2Core_pixelsOut_payload_pixel;
  wire                rChannelPart2Core_pixelsOut_payload_frameStart;
  wire                rChannelPart2Core_pixelsOut_payload_rowEnd;
  wire                rChannelPart2Core_pixelsOut_payload_inpValid;
  wire                rChannelPart2Core_startOut;
  wire                rChannelPart2Core_inpTwoDoneOut;
  wire                rChannelPart3Core_pixelsIn_ready;
  wire                rChannelPart3Core_pixelsOut_valid;
  wire       [7:0]    rChannelPart3Core_pixelsOut_payload_pixel;
  wire                rChannelPart3Core_pixelsOut_payload_frameStart;
  wire                rChannelPart3Core_pixelsOut_payload_rowEnd;
  wire                rChannelPart3Core_inpThreeDoneOut;
  wire                channelCombiner_bPixelChannelIn_ready;
  wire                channelCombiner_gPixelChannelIn_ready;
  wire                channelCombiner_rPixelChannelIn_ready;
  wire                channelCombiner_allPixelChannelOut_valid;
  wire       [31:0]   channelCombiner_allPixelChannelOut_payload_pixel;
  wire                channelCombiner_allPixelChannelOut_payload_frameStart;
  wire                channelCombiner_allPixelChannelOut_payload_rowEnd;
  wire                inpConfig_1_axiLiteSignal_aw_ready;
  wire                inpConfig_1_axiLiteSignal_w_ready;
  wire                inpConfig_1_axiLiteSignal_b_valid;
  wire       [1:0]    inpConfig_1_axiLiteSignal_b_payload_resp;
  wire                inpConfig_1_axiLiteSignal_ar_ready;
  wire                inpConfig_1_axiLiteSignal_r_valid;
  wire       [31:0]   inpConfig_1_axiLiteSignal_r_payload_data;
  wire       [1:0]    inpConfig_1_axiLiteSignal_r_payload_resp;
  wire       [9:0]    inpConfig_1_srcWidth;
  wire       [9:0]    inpConfig_1_srcHeight;
  wire       [7:0]    inpConfig_1_threshold;
  wire                inpConfig_1_apStart;
  reg                 rDone;
  reg                 gDone;
  reg                 bDone;
  wire                allChannelDone;

  DDRDataWrapper ddrDataWrapper_1 (
    .ddrIn_valid                  (ddrDataIn_valid                               ), //i
    .ddrIn_ready                  (ddrDataWrapper_1_ddrIn_ready                  ), //o
    .ddrIn_payload                (ddrDataIn_payload[31:0]                       ), //i
    .pixelsOut_valid              (ddrDataWrapper_1_pixelsOut_valid              ), //o
    .pixelsOut_ready              (channelDispatcher_allPixelChannelIn_ready     ), //i
    .pixelsOut_payload_pixel      (ddrDataWrapper_1_pixelsOut_payload_pixel[31:0]), //o
    .pixelsOut_payload_frameStart (ddrDataWrapper_1_pixelsOut_payload_frameStart ), //o
    .pixelsOut_payload_rowEnd     (ddrDataWrapper_1_pixelsOut_payload_rowEnd     ), //o
    .inpDone                      (allChannelDone                                ), //i
    .bmpWidth                     (inpConfig_1_srcWidth[9:0]                     ), //i
    .clk                          (clk                                           ), //i
    .resetn                       (resetn                                        )  //i
  );
  ChannelMasterTransformer channelDispatcher (
    .allPixelChannelIn_valid              (ddrDataWrapper_1_pixelsOut_valid                     ), //i
    .allPixelChannelIn_ready              (channelDispatcher_allPixelChannelIn_ready            ), //o
    .allPixelChannelIn_payload_pixel      (ddrDataWrapper_1_pixelsOut_payload_pixel[31:0]       ), //i
    .allPixelChannelIn_payload_frameStart (ddrDataWrapper_1_pixelsOut_payload_frameStart        ), //i
    .allPixelChannelIn_payload_rowEnd     (ddrDataWrapper_1_pixelsOut_payload_rowEnd            ), //i
    .bPixelChannelOut_valid               (channelDispatcher_bPixelChannelOut_valid             ), //o
    .bPixelChannelOut_ready               (bChannelPart1Core_pixelsIn_ready                     ), //i
    .bPixelChannelOut_payload_pixel       (channelDispatcher_bPixelChannelOut_payload_pixel[7:0]), //o
    .bPixelChannelOut_payload_frameStart  (channelDispatcher_bPixelChannelOut_payload_frameStart), //o
    .bPixelChannelOut_payload_rowEnd      (channelDispatcher_bPixelChannelOut_payload_rowEnd    ), //o
    .gPixelChannelOut_valid               (channelDispatcher_gPixelChannelOut_valid             ), //o
    .gPixelChannelOut_ready               (gChannelPart1Core_pixelsIn_ready                     ), //i
    .gPixelChannelOut_payload_pixel       (channelDispatcher_gPixelChannelOut_payload_pixel[7:0]), //o
    .gPixelChannelOut_payload_frameStart  (channelDispatcher_gPixelChannelOut_payload_frameStart), //o
    .gPixelChannelOut_payload_rowEnd      (channelDispatcher_gPixelChannelOut_payload_rowEnd    ), //o
    .rPixelChannelOut_valid               (channelDispatcher_rPixelChannelOut_valid             ), //o
    .rPixelChannelOut_ready               (rChannelPart1Core_pixelsIn_ready                     ), //i
    .rPixelChannelOut_payload_pixel       (channelDispatcher_rPixelChannelOut_payload_pixel[7:0]), //o
    .rPixelChannelOut_payload_frameStart  (channelDispatcher_rPixelChannelOut_payload_frameStart), //o
    .rPixelChannelOut_payload_rowEnd      (channelDispatcher_rPixelChannelOut_payload_rowEnd    ), //o
    .clk                                  (clk                                                  ), //i
    .resetn                               (resetn                                               )  //i
  );
  SuperResolutionPart1 bChannelPart1Core (
    .pixelsIn_valid               (channelDispatcher_bPixelChannelOut_valid             ), //i
    .pixelsIn_ready               (bChannelPart1Core_pixelsIn_ready                     ), //o
    .pixelsIn_payload_pixel       (channelDispatcher_bPixelChannelOut_payload_pixel[7:0]), //i
    .pixelsIn_payload_frameStart  (channelDispatcher_bPixelChannelOut_payload_frameStart), //i
    .pixelsIn_payload_rowEnd      (channelDispatcher_bPixelChannelOut_payload_rowEnd    ), //i
    .startIn                      (inpConfig_1_apStart                                  ), //i
    .inpTwoDoneIn                 (bChannelPart2Core_inpTwoDoneOut                      ), //i
    .inpThreeDoneIn               (bChannelPart3Core_inpThreeDoneOut                    ), //i
    .pixelsOut_valid              (bChannelPart1Core_pixelsOut_valid                    ), //o
    .pixelsOut_ready              (bChannelPart2Core_pixelsIn_ready                     ), //i
    .pixelsOut_payload_pixel      (bChannelPart1Core_pixelsOut_payload_pixel[7:0]       ), //o
    .pixelsOut_payload_frameStart (bChannelPart1Core_pixelsOut_payload_frameStart       ), //o
    .pixelsOut_payload_rowEnd     (bChannelPart1Core_pixelsOut_payload_rowEnd           ), //o
    .startOut                     (bChannelPart1Core_startOut                           ), //o
    .inpDoneOut                   (bChannelPart1Core_inpDoneOut                         ), //o
    .thresholdIn                  (inpConfig_1_threshold[7:0]                           ), //i
    .widthIn                      (inpConfig_1_srcWidth[9:0]                            ), //i
    .heightIn                     (inpConfig_1_srcHeight[9:0]                           ), //i
    .clk                          (clk                                                  ), //i
    .resetn                       (resetn                                               )  //i
  );
  SuperResolutionPart2 bChannelPart2Core (
    .pixelsIn_valid               (bChannelPart1Core_pixelsOut_valid             ), //i
    .pixelsIn_ready               (bChannelPart2Core_pixelsIn_ready              ), //o
    .pixelsIn_payload_pixel       (bChannelPart1Core_pixelsOut_payload_pixel[7:0]), //i
    .pixelsIn_payload_frameStart  (bChannelPart1Core_pixelsOut_payload_frameStart), //i
    .pixelsIn_payload_rowEnd      (bChannelPart1Core_pixelsOut_payload_rowEnd    ), //i
    .startIn                      (bChannelPart1Core_startOut                    ), //i
    .inpThreeDoneIn               (bChannelPart3Core_inpThreeDoneOut             ), //i
    .pixelsOut_valid              (bChannelPart2Core_pixelsOut_valid             ), //o
    .pixelsOut_ready              (bChannelPart3Core_pixelsIn_ready              ), //i
    .pixelsOut_payload_pixel      (bChannelPart2Core_pixelsOut_payload_pixel[7:0]), //o
    .pixelsOut_payload_frameStart (bChannelPart2Core_pixelsOut_payload_frameStart), //o
    .pixelsOut_payload_rowEnd     (bChannelPart2Core_pixelsOut_payload_rowEnd    ), //o
    .pixelsOut_payload_inpValid   (bChannelPart2Core_pixelsOut_payload_inpValid  ), //o
    .startOut                     (bChannelPart2Core_startOut                    ), //o
    .inpTwoDoneOut                (bChannelPart2Core_inpTwoDoneOut               ), //o
    .thresholdIn                  (inpConfig_1_threshold[7:0]                    ), //i
    .widthIn                      (inpConfig_1_srcWidth[9:0]                     ), //i
    .heightIn                     (inpConfig_1_srcHeight[9:0]                    ), //i
    .clk                          (clk                                           ), //i
    .resetn                       (resetn                                        )  //i
  );
  SuperResolutionPart3 bChannelPart3Core (
    .pixelsIn_valid               (bChannelPart2Core_pixelsOut_valid             ), //i
    .pixelsIn_ready               (bChannelPart3Core_pixelsIn_ready              ), //o
    .pixelsIn_payload_pixel       (bChannelPart2Core_pixelsOut_payload_pixel[7:0]), //i
    .pixelsIn_payload_frameStart  (bChannelPart2Core_pixelsOut_payload_frameStart), //i
    .pixelsIn_payload_rowEnd      (bChannelPart2Core_pixelsOut_payload_rowEnd    ), //i
    .pixelsIn_payload_inpValid    (bChannelPart2Core_pixelsOut_payload_inpValid  ), //i
    .startIn                      (bChannelPart2Core_startOut                    ), //i
    .pixelsOut_valid              (bChannelPart3Core_pixelsOut_valid             ), //o
    .pixelsOut_ready              (channelCombiner_bPixelChannelIn_ready         ), //i
    .pixelsOut_payload_pixel      (bChannelPart3Core_pixelsOut_payload_pixel[7:0]), //o
    .pixelsOut_payload_frameStart (bChannelPart3Core_pixelsOut_payload_frameStart), //o
    .pixelsOut_payload_rowEnd     (bChannelPart3Core_pixelsOut_payload_rowEnd    ), //o
    .inpThreeDoneOut              (bChannelPart3Core_inpThreeDoneOut             ), //o
    .thresholdIn                  (inpConfig_1_threshold[7:0]                    ), //i
    .widthIn                      (inpConfig_1_srcWidth[9:0]                     ), //i
    .heightIn                     (inpConfig_1_srcHeight[9:0]                    ), //i
    .clk                          (clk                                           ), //i
    .resetn                       (resetn                                        )  //i
  );
  SuperResolutionPart1_1 gChannelPart1Core (
    .pixelsIn_valid               (channelDispatcher_gPixelChannelOut_valid             ), //i
    .pixelsIn_ready               (gChannelPart1Core_pixelsIn_ready                     ), //o
    .pixelsIn_payload_pixel       (channelDispatcher_gPixelChannelOut_payload_pixel[7:0]), //i
    .pixelsIn_payload_frameStart  (channelDispatcher_gPixelChannelOut_payload_frameStart), //i
    .pixelsIn_payload_rowEnd      (channelDispatcher_gPixelChannelOut_payload_rowEnd    ), //i
    .startIn                      (inpConfig_1_apStart                                  ), //i
    .inpTwoDoneIn                 (gChannelPart2Core_inpTwoDoneOut                      ), //i
    .inpThreeDoneIn               (gChannelPart3Core_inpThreeDoneOut                    ), //i
    .pixelsOut_valid              (gChannelPart1Core_pixelsOut_valid                    ), //o
    .pixelsOut_ready              (gChannelPart2Core_pixelsIn_ready                     ), //i
    .pixelsOut_payload_pixel      (gChannelPart1Core_pixelsOut_payload_pixel[7:0]       ), //o
    .pixelsOut_payload_frameStart (gChannelPart1Core_pixelsOut_payload_frameStart       ), //o
    .pixelsOut_payload_rowEnd     (gChannelPart1Core_pixelsOut_payload_rowEnd           ), //o
    .startOut                     (gChannelPart1Core_startOut                           ), //o
    .inpDoneOut                   (gChannelPart1Core_inpDoneOut                         ), //o
    .thresholdIn                  (inpConfig_1_threshold[7:0]                           ), //i
    .widthIn                      (inpConfig_1_srcWidth[9:0]                            ), //i
    .heightIn                     (inpConfig_1_srcHeight[9:0]                           ), //i
    .clk                          (clk                                                  ), //i
    .resetn                       (resetn                                               )  //i
  );
  SuperResolutionPart2_1 gChannelPart2Core (
    .pixelsIn_valid               (gChannelPart1Core_pixelsOut_valid             ), //i
    .pixelsIn_ready               (gChannelPart2Core_pixelsIn_ready              ), //o
    .pixelsIn_payload_pixel       (gChannelPart1Core_pixelsOut_payload_pixel[7:0]), //i
    .pixelsIn_payload_frameStart  (gChannelPart1Core_pixelsOut_payload_frameStart), //i
    .pixelsIn_payload_rowEnd      (gChannelPart1Core_pixelsOut_payload_rowEnd    ), //i
    .startIn                      (gChannelPart1Core_startOut                    ), //i
    .inpThreeDoneIn               (gChannelPart3Core_inpThreeDoneOut             ), //i
    .pixelsOut_valid              (gChannelPart2Core_pixelsOut_valid             ), //o
    .pixelsOut_ready              (gChannelPart3Core_pixelsIn_ready              ), //i
    .pixelsOut_payload_pixel      (gChannelPart2Core_pixelsOut_payload_pixel[7:0]), //o
    .pixelsOut_payload_frameStart (gChannelPart2Core_pixelsOut_payload_frameStart), //o
    .pixelsOut_payload_rowEnd     (gChannelPart2Core_pixelsOut_payload_rowEnd    ), //o
    .pixelsOut_payload_inpValid   (gChannelPart2Core_pixelsOut_payload_inpValid  ), //o
    .startOut                     (gChannelPart2Core_startOut                    ), //o
    .inpTwoDoneOut                (gChannelPart2Core_inpTwoDoneOut               ), //o
    .thresholdIn                  (inpConfig_1_threshold[7:0]                    ), //i
    .widthIn                      (inpConfig_1_srcWidth[9:0]                     ), //i
    .heightIn                     (inpConfig_1_srcHeight[9:0]                    ), //i
    .clk                          (clk                                           ), //i
    .resetn                       (resetn                                        )  //i
  );
  SuperResolutionPart3_1 gChannelPart3Core (
    .pixelsIn_valid               (gChannelPart2Core_pixelsOut_valid             ), //i
    .pixelsIn_ready               (gChannelPart3Core_pixelsIn_ready              ), //o
    .pixelsIn_payload_pixel       (gChannelPart2Core_pixelsOut_payload_pixel[7:0]), //i
    .pixelsIn_payload_frameStart  (gChannelPart2Core_pixelsOut_payload_frameStart), //i
    .pixelsIn_payload_rowEnd      (gChannelPart2Core_pixelsOut_payload_rowEnd    ), //i
    .pixelsIn_payload_inpValid    (gChannelPart2Core_pixelsOut_payload_inpValid  ), //i
    .startIn                      (gChannelPart2Core_startOut                    ), //i
    .pixelsOut_valid              (gChannelPart3Core_pixelsOut_valid             ), //o
    .pixelsOut_ready              (channelCombiner_gPixelChannelIn_ready         ), //i
    .pixelsOut_payload_pixel      (gChannelPart3Core_pixelsOut_payload_pixel[7:0]), //o
    .pixelsOut_payload_frameStart (gChannelPart3Core_pixelsOut_payload_frameStart), //o
    .pixelsOut_payload_rowEnd     (gChannelPart3Core_pixelsOut_payload_rowEnd    ), //o
    .inpThreeDoneOut              (gChannelPart3Core_inpThreeDoneOut             ), //o
    .thresholdIn                  (inpConfig_1_threshold[7:0]                    ), //i
    .widthIn                      (inpConfig_1_srcWidth[9:0]                     ), //i
    .heightIn                     (inpConfig_1_srcHeight[9:0]                    ), //i
    .clk                          (clk                                           ), //i
    .resetn                       (resetn                                        )  //i
  );
  SuperResolutionPart1_2 rChannelPart1Core (
    .pixelsIn_valid               (channelDispatcher_rPixelChannelOut_valid             ), //i
    .pixelsIn_ready               (rChannelPart1Core_pixelsIn_ready                     ), //o
    .pixelsIn_payload_pixel       (channelDispatcher_rPixelChannelOut_payload_pixel[7:0]), //i
    .pixelsIn_payload_frameStart  (channelDispatcher_rPixelChannelOut_payload_frameStart), //i
    .pixelsIn_payload_rowEnd      (channelDispatcher_rPixelChannelOut_payload_rowEnd    ), //i
    .startIn                      (inpConfig_1_apStart                                  ), //i
    .inpTwoDoneIn                 (rChannelPart2Core_inpTwoDoneOut                      ), //i
    .inpThreeDoneIn               (rChannelPart3Core_inpThreeDoneOut                    ), //i
    .pixelsOut_valid              (rChannelPart1Core_pixelsOut_valid                    ), //o
    .pixelsOut_ready              (rChannelPart2Core_pixelsIn_ready                     ), //i
    .pixelsOut_payload_pixel      (rChannelPart1Core_pixelsOut_payload_pixel[7:0]       ), //o
    .pixelsOut_payload_frameStart (rChannelPart1Core_pixelsOut_payload_frameStart       ), //o
    .pixelsOut_payload_rowEnd     (rChannelPart1Core_pixelsOut_payload_rowEnd           ), //o
    .startOut                     (rChannelPart1Core_startOut                           ), //o
    .inpDoneOut                   (rChannelPart1Core_inpDoneOut                         ), //o
    .thresholdIn                  (inpConfig_1_threshold[7:0]                           ), //i
    .widthIn                      (inpConfig_1_srcWidth[9:0]                            ), //i
    .heightIn                     (inpConfig_1_srcHeight[9:0]                           ), //i
    .clk                          (clk                                                  ), //i
    .resetn                       (resetn                                               )  //i
  );
  SuperResolutionPart2_2 rChannelPart2Core (
    .pixelsIn_valid               (rChannelPart1Core_pixelsOut_valid             ), //i
    .pixelsIn_ready               (rChannelPart2Core_pixelsIn_ready              ), //o
    .pixelsIn_payload_pixel       (rChannelPart1Core_pixelsOut_payload_pixel[7:0]), //i
    .pixelsIn_payload_frameStart  (rChannelPart1Core_pixelsOut_payload_frameStart), //i
    .pixelsIn_payload_rowEnd      (rChannelPart1Core_pixelsOut_payload_rowEnd    ), //i
    .startIn                      (rChannelPart1Core_startOut                    ), //i
    .inpThreeDoneIn               (rChannelPart3Core_inpThreeDoneOut             ), //i
    .pixelsOut_valid              (rChannelPart2Core_pixelsOut_valid             ), //o
    .pixelsOut_ready              (rChannelPart3Core_pixelsIn_ready              ), //i
    .pixelsOut_payload_pixel      (rChannelPart2Core_pixelsOut_payload_pixel[7:0]), //o
    .pixelsOut_payload_frameStart (rChannelPart2Core_pixelsOut_payload_frameStart), //o
    .pixelsOut_payload_rowEnd     (rChannelPart2Core_pixelsOut_payload_rowEnd    ), //o
    .pixelsOut_payload_inpValid   (rChannelPart2Core_pixelsOut_payload_inpValid  ), //o
    .startOut                     (rChannelPart2Core_startOut                    ), //o
    .inpTwoDoneOut                (rChannelPart2Core_inpTwoDoneOut               ), //o
    .thresholdIn                  (inpConfig_1_threshold[7:0]                    ), //i
    .widthIn                      (inpConfig_1_srcWidth[9:0]                     ), //i
    .heightIn                     (inpConfig_1_srcHeight[9:0]                    ), //i
    .clk                          (clk                                           ), //i
    .resetn                       (resetn                                        )  //i
  );
  SuperResolutionPart3_2 rChannelPart3Core (
    .pixelsIn_valid               (rChannelPart2Core_pixelsOut_valid             ), //i
    .pixelsIn_ready               (rChannelPart3Core_pixelsIn_ready              ), //o
    .pixelsIn_payload_pixel       (rChannelPart2Core_pixelsOut_payload_pixel[7:0]), //i
    .pixelsIn_payload_frameStart  (rChannelPart2Core_pixelsOut_payload_frameStart), //i
    .pixelsIn_payload_rowEnd      (rChannelPart2Core_pixelsOut_payload_rowEnd    ), //i
    .pixelsIn_payload_inpValid    (rChannelPart2Core_pixelsOut_payload_inpValid  ), //i
    .startIn                      (rChannelPart2Core_startOut                    ), //i
    .pixelsOut_valid              (rChannelPart3Core_pixelsOut_valid             ), //o
    .pixelsOut_ready              (channelCombiner_rPixelChannelIn_ready         ), //i
    .pixelsOut_payload_pixel      (rChannelPart3Core_pixelsOut_payload_pixel[7:0]), //o
    .pixelsOut_payload_frameStart (rChannelPart3Core_pixelsOut_payload_frameStart), //o
    .pixelsOut_payload_rowEnd     (rChannelPart3Core_pixelsOut_payload_rowEnd    ), //o
    .inpThreeDoneOut              (rChannelPart3Core_inpThreeDoneOut             ), //o
    .thresholdIn                  (inpConfig_1_threshold[7:0]                    ), //i
    .widthIn                      (inpConfig_1_srcWidth[9:0]                     ), //i
    .heightIn                     (inpConfig_1_srcHeight[9:0]                    ), //i
    .clk                          (clk                                           ), //i
    .resetn                       (resetn                                        )  //i
  );
  ChannelSlaveTransformer channelCombiner (
    .bPixelChannelIn_valid                 (bChannelPart3Core_pixelsOut_valid                     ), //i
    .bPixelChannelIn_ready                 (channelCombiner_bPixelChannelIn_ready                 ), //o
    .bPixelChannelIn_payload_pixel         (bChannelPart3Core_pixelsOut_payload_pixel[7:0]        ), //i
    .bPixelChannelIn_payload_frameStart    (bChannelPart3Core_pixelsOut_payload_frameStart        ), //i
    .bPixelChannelIn_payload_rowEnd        (bChannelPart3Core_pixelsOut_payload_rowEnd            ), //i
    .gPixelChannelIn_valid                 (gChannelPart3Core_pixelsOut_valid                     ), //i
    .gPixelChannelIn_ready                 (channelCombiner_gPixelChannelIn_ready                 ), //o
    .gPixelChannelIn_payload_pixel         (gChannelPart3Core_pixelsOut_payload_pixel[7:0]        ), //i
    .gPixelChannelIn_payload_frameStart    (gChannelPart3Core_pixelsOut_payload_frameStart        ), //i
    .gPixelChannelIn_payload_rowEnd        (gChannelPart3Core_pixelsOut_payload_rowEnd            ), //i
    .rPixelChannelIn_valid                 (rChannelPart3Core_pixelsOut_valid                     ), //i
    .rPixelChannelIn_ready                 (channelCombiner_rPixelChannelIn_ready                 ), //o
    .rPixelChannelIn_payload_pixel         (rChannelPart3Core_pixelsOut_payload_pixel[7:0]        ), //i
    .rPixelChannelIn_payload_frameStart    (rChannelPart3Core_pixelsOut_payload_frameStart        ), //i
    .rPixelChannelIn_payload_rowEnd        (rChannelPart3Core_pixelsOut_payload_rowEnd            ), //i
    .allPixelChannelOut_valid              (channelCombiner_allPixelChannelOut_valid              ), //o
    .allPixelChannelOut_ready              (inpDataOut_ready                                      ), //i
    .allPixelChannelOut_payload_pixel      (channelCombiner_allPixelChannelOut_payload_pixel[31:0]), //o
    .allPixelChannelOut_payload_frameStart (channelCombiner_allPixelChannelOut_payload_frameStart ), //o
    .allPixelChannelOut_payload_rowEnd     (channelCombiner_allPixelChannelOut_payload_rowEnd     ), //o
    .clk                                   (clk                                                   ), //i
    .resetn                                (resetn                                                )  //i
  );
  InpConfig inpConfig_1 (
    .axiLiteSignal_aw_valid        (ipConfig_aw_valid                             ), //i
    .axiLiteSignal_aw_ready        (inpConfig_1_axiLiteSignal_aw_ready            ), //o
    .axiLiteSignal_aw_payload_addr (ipConfig_aw_payload_addr[31:0]                ), //i
    .axiLiteSignal_aw_payload_prot (ipConfig_aw_payload_prot[2:0]                 ), //i
    .axiLiteSignal_w_valid         (ipConfig_w_valid                              ), //i
    .axiLiteSignal_w_ready         (inpConfig_1_axiLiteSignal_w_ready             ), //o
    .axiLiteSignal_w_payload_data  (ipConfig_w_payload_data[31:0]                 ), //i
    .axiLiteSignal_w_payload_strb  (ipConfig_w_payload_strb[3:0]                  ), //i
    .axiLiteSignal_b_valid         (inpConfig_1_axiLiteSignal_b_valid             ), //o
    .axiLiteSignal_b_ready         (ipConfig_b_ready                              ), //i
    .axiLiteSignal_b_payload_resp  (inpConfig_1_axiLiteSignal_b_payload_resp[1:0] ), //o
    .axiLiteSignal_ar_valid        (ipConfig_ar_valid                             ), //i
    .axiLiteSignal_ar_ready        (inpConfig_1_axiLiteSignal_ar_ready            ), //o
    .axiLiteSignal_ar_payload_addr (ipConfig_ar_payload_addr[31:0]                ), //i
    .axiLiteSignal_ar_payload_prot (ipConfig_ar_payload_prot[2:0]                 ), //i
    .axiLiteSignal_r_valid         (inpConfig_1_axiLiteSignal_r_valid             ), //o
    .axiLiteSignal_r_ready         (ipConfig_r_ready                              ), //i
    .axiLiteSignal_r_payload_data  (inpConfig_1_axiLiteSignal_r_payload_data[31:0]), //o
    .axiLiteSignal_r_payload_resp  (inpConfig_1_axiLiteSignal_r_payload_resp[1:0] ), //o
    .apDone                        (allChannelDone                                ), //i
    .srcWidth                      (inpConfig_1_srcWidth[9:0]                     ), //o
    .srcHeight                     (inpConfig_1_srcHeight[9:0]                    ), //o
    .threshold                     (inpConfig_1_threshold[7:0]                    ), //o
    .apStart                       (inpConfig_1_apStart                           ), //o
    .clk                           (clk                                           ), //i
    .resetn                        (resetn                                        )  //i
  );
  assign allChannelDone = ((rDone && gDone) && bDone);
  assign ddrDataIn_ready = ddrDataWrapper_1_ddrIn_ready;
  assign ipConfig_aw_ready = inpConfig_1_axiLiteSignal_aw_ready;
  assign ipConfig_w_ready = inpConfig_1_axiLiteSignal_w_ready;
  assign ipConfig_b_valid = inpConfig_1_axiLiteSignal_b_valid;
  assign ipConfig_b_payload_resp = inpConfig_1_axiLiteSignal_b_payload_resp;
  assign ipConfig_ar_ready = inpConfig_1_axiLiteSignal_ar_ready;
  assign ipConfig_r_valid = inpConfig_1_axiLiteSignal_r_valid;
  assign ipConfig_r_payload_data = inpConfig_1_axiLiteSignal_r_payload_data;
  assign ipConfig_r_payload_resp = inpConfig_1_axiLiteSignal_r_payload_resp;
  assign inpDataOut_valid = channelCombiner_allPixelChannelOut_valid;
  assign inpDataOut_payload_pixel = channelCombiner_allPixelChannelOut_payload_pixel;
  assign inpDataOut_payload_frameStart = channelCombiner_allPixelChannelOut_payload_frameStart;
  assign inpDataOut_payload_rowEnd = channelCombiner_allPixelChannelOut_payload_rowEnd;
  always @(posedge clk or negedge resetn) begin
    if(!resetn) begin
      rDone <= 1'b0;
      gDone <= 1'b0;
      bDone <= 1'b0;
    end else begin
      rDone <= rChannelPart1Core_inpDoneOut;
      gDone <= gChannelPart1Core_inpDoneOut;
      bDone <= bChannelPart1Core_inpDoneOut;
      if(allChannelDone) begin
        rDone <= 1'b0;
        gDone <= 1'b0;
        bDone <= 1'b0;
      end
    end
  end


endmodule

module InpConfig (
  input               axiLiteSignal_aw_valid,
  output              axiLiteSignal_aw_ready,
  input      [31:0]   axiLiteSignal_aw_payload_addr,
  input      [2:0]    axiLiteSignal_aw_payload_prot,
  input               axiLiteSignal_w_valid,
  output              axiLiteSignal_w_ready,
  input      [31:0]   axiLiteSignal_w_payload_data,
  input      [3:0]    axiLiteSignal_w_payload_strb,
  output              axiLiteSignal_b_valid,
  input               axiLiteSignal_b_ready,
  output     [1:0]    axiLiteSignal_b_payload_resp,
  input               axiLiteSignal_ar_valid,
  output              axiLiteSignal_ar_ready,
  input      [31:0]   axiLiteSignal_ar_payload_addr,
  input      [2:0]    axiLiteSignal_ar_payload_prot,
  output reg          axiLiteSignal_r_valid,
  input               axiLiteSignal_r_ready,
  output reg [31:0]   axiLiteSignal_r_payload_data,
  output     [1:0]    axiLiteSignal_r_payload_resp,
  input               apDone,
  output     [9:0]    srcWidth,
  output     [9:0]    srcHeight,
  output     [7:0]    threshold,
  output              apStart,
  input               clk,
  input               resetn
);

  wire       [9:0]    CICC1851_axiLiteSignal_r_payload_data;
  wire       [9:0]    CICC1851_axiLiteSignal_r_payload_data_1;
  wire       [7:0]    CICC1851_axiLiteSignal_r_payload_data_2;
  wire       [0:0]    CICC1851_axiLiteSignal_r_payload_data_3;
  reg        [9:0]    regSrcW;
  reg        [9:0]    regSrcH;
  reg        [7:0]    regThreshold;
  reg                 regApStart;
  reg        [7:0]    regWrAddr;
  reg        [7:0]    regRAddr;
  reg                 updateWrAddr;
  reg                 updateRAddr;
  reg                 writeSuccess;
  wire                axiLiteSignal_aw_fire;
  wire                axiLiteSignal_aw_fire_1;
  wire                axiLiteSignal_w_fire;
  wire                axiLiteSignal_w_fire_1;
  wire                axiLiteSignal_w_fire_2;
  wire                axiLiteSignal_b_fire;
  wire                axiLiteSignal_ar_fire;
  wire                axiLiteSignal_ar_fire_1;
  wire                axiLiteSignal_r_fire;
  wire                when_InpConfig_l69;

  assign CICC1851_axiLiteSignal_r_payload_data = regSrcW;
  assign CICC1851_axiLiteSignal_r_payload_data_1 = regSrcH;
  assign CICC1851_axiLiteSignal_r_payload_data_2 = regThreshold;
  assign CICC1851_axiLiteSignal_r_payload_data_3 = regApStart;
  assign axiLiteSignal_aw_ready = updateWrAddr;
  assign axiLiteSignal_aw_fire = (axiLiteSignal_aw_valid && axiLiteSignal_aw_ready);
  assign axiLiteSignal_aw_fire_1 = (axiLiteSignal_aw_valid && axiLiteSignal_aw_ready);
  assign axiLiteSignal_w_fire = (axiLiteSignal_w_valid && axiLiteSignal_w_ready);
  assign axiLiteSignal_w_ready = (! updateWrAddr);
  assign axiLiteSignal_w_fire_1 = (axiLiteSignal_w_valid && axiLiteSignal_w_ready);
  assign axiLiteSignal_w_fire_2 = (axiLiteSignal_w_valid && axiLiteSignal_w_ready);
  assign axiLiteSignal_b_fire = (axiLiteSignal_b_valid && axiLiteSignal_b_ready);
  assign axiLiteSignal_b_valid = writeSuccess;
  assign axiLiteSignal_b_payload_resp = 2'b00;
  assign axiLiteSignal_ar_ready = updateRAddr;
  assign axiLiteSignal_ar_fire = (axiLiteSignal_ar_valid && axiLiteSignal_ar_ready);
  assign axiLiteSignal_ar_fire_1 = (axiLiteSignal_ar_valid && axiLiteSignal_ar_ready);
  assign axiLiteSignal_r_fire = (axiLiteSignal_r_valid && axiLiteSignal_r_ready);
  assign axiLiteSignal_r_payload_resp = 2'b00;
  assign when_InpConfig_l69 = (! updateRAddr);
  always @(*) begin
    if(when_InpConfig_l69) begin
      axiLiteSignal_r_valid = 1'b1;
    end else begin
      axiLiteSignal_r_valid = 1'b1;
    end
  end

  always @(*) begin
    if(when_InpConfig_l69) begin
      case(regRAddr)
        8'h04 : begin
          axiLiteSignal_r_payload_data = {22'd0, CICC1851_axiLiteSignal_r_payload_data};
        end
        8'h08 : begin
          axiLiteSignal_r_payload_data = {22'd0, CICC1851_axiLiteSignal_r_payload_data_1};
        end
        8'h0c : begin
          axiLiteSignal_r_payload_data = {24'd0, CICC1851_axiLiteSignal_r_payload_data_2};
        end
        8'h10 : begin
          axiLiteSignal_r_payload_data = {31'd0, CICC1851_axiLiteSignal_r_payload_data_3};
        end
        default : begin
          axiLiteSignal_r_payload_data = 32'h0;
        end
      endcase
    end else begin
      axiLiteSignal_r_payload_data = 32'h0;
    end
  end

  assign srcWidth = regSrcW;
  assign srcHeight = regSrcH;
  assign threshold = regThreshold;
  assign apStart = regApStart;
  always @(posedge clk or negedge resetn) begin
    if(!resetn) begin
      regSrcW <= 10'h0;
      regSrcH <= 10'h0;
      regThreshold <= 8'hff;
      regApStart <= 1'b0;
      regWrAddr <= 8'hff;
      regRAddr <= 8'hff;
      updateWrAddr <= 1'b1;
      updateRAddr <= 1'b1;
      writeSuccess <= 1'b0;
    end else begin
      if(axiLiteSignal_aw_fire) begin
        regWrAddr <= axiLiteSignal_aw_payload_addr[7 : 0];
      end
      if(axiLiteSignal_aw_fire_1) begin
        updateWrAddr <= 1'b0;
      end else begin
        if(axiLiteSignal_w_fire) begin
          updateWrAddr <= 1'b1;
        end
      end
      if(axiLiteSignal_w_fire_1) begin
        case(regWrAddr)
          8'h04 : begin
            regSrcW <= axiLiteSignal_w_payload_data[9 : 0];
          end
          8'h08 : begin
            regSrcH <= axiLiteSignal_w_payload_data[9 : 0];
          end
          8'h0c : begin
            regThreshold <= axiLiteSignal_w_payload_data[7 : 0];
          end
          8'h10 : begin
            regApStart <= axiLiteSignal_w_payload_data[0];
          end
          default : begin
          end
        endcase
      end
      if(axiLiteSignal_w_fire_2) begin
        writeSuccess <= 1'b1;
      end else begin
        if(axiLiteSignal_b_fire) begin
          writeSuccess <= 1'b0;
        end
      end
      if(axiLiteSignal_ar_fire) begin
        regRAddr <= axiLiteSignal_ar_payload_addr[7 : 0];
      end
      if(axiLiteSignal_ar_fire_1) begin
        updateRAddr <= 1'b0;
      end else begin
        if(axiLiteSignal_r_fire) begin
          updateRAddr <= 1'b1;
        end
      end
      if(apDone) begin
        regApStart <= 1'b0;
      end
    end
  end


endmodule

module ChannelSlaveTransformer (
  input               bPixelChannelIn_valid,
  output reg          bPixelChannelIn_ready,
  input      [7:0]    bPixelChannelIn_payload_pixel,
  input               bPixelChannelIn_payload_frameStart,
  input               bPixelChannelIn_payload_rowEnd,
  input               gPixelChannelIn_valid,
  output reg          gPixelChannelIn_ready,
  input      [7:0]    gPixelChannelIn_payload_pixel,
  input               gPixelChannelIn_payload_frameStart,
  input               gPixelChannelIn_payload_rowEnd,
  input               rPixelChannelIn_valid,
  output reg          rPixelChannelIn_ready,
  input      [7:0]    rPixelChannelIn_payload_pixel,
  input               rPixelChannelIn_payload_frameStart,
  input               rPixelChannelIn_payload_rowEnd,
  output              allPixelChannelOut_valid,
  input               allPixelChannelOut_ready,
  output     [31:0]   allPixelChannelOut_payload_pixel,
  output              allPixelChannelOut_payload_frameStart,
  output              allPixelChannelOut_payload_rowEnd,
  input               clk,
  input               resetn
);

  wire                bPixelChannelIn_m2sPipe_valid;
  wire                bPixelChannelIn_m2sPipe_ready;
  wire       [7:0]    bPixelChannelIn_m2sPipe_payload_pixel;
  wire                bPixelChannelIn_m2sPipe_payload_frameStart;
  wire                bPixelChannelIn_m2sPipe_payload_rowEnd;
  reg                 bPixelChannelIn_rValid;
  reg        [7:0]    bPixelChannelIn_rData_pixel;
  reg                 bPixelChannelIn_rData_frameStart;
  reg                 bPixelChannelIn_rData_rowEnd;
  wire                when_Stream_l368;
  wire                gPixelChannelIn_m2sPipe_valid;
  wire                gPixelChannelIn_m2sPipe_ready;
  wire       [7:0]    gPixelChannelIn_m2sPipe_payload_pixel;
  wire                gPixelChannelIn_m2sPipe_payload_frameStart;
  wire                gPixelChannelIn_m2sPipe_payload_rowEnd;
  reg                 gPixelChannelIn_rValid;
  reg        [7:0]    gPixelChannelIn_rData_pixel;
  reg                 gPixelChannelIn_rData_frameStart;
  reg                 gPixelChannelIn_rData_rowEnd;
  wire                when_Stream_l368_1;
  wire                rPixelChannelIn_m2sPipe_valid;
  wire                rPixelChannelIn_m2sPipe_ready;
  wire       [7:0]    rPixelChannelIn_m2sPipe_payload_pixel;
  wire                rPixelChannelIn_m2sPipe_payload_frameStart;
  wire                rPixelChannelIn_m2sPipe_payload_rowEnd;
  reg                 rPixelChannelIn_rValid;
  reg        [7:0]    rPixelChannelIn_rData_pixel;
  reg                 rPixelChannelIn_rData_frameStart;
  reg                 rPixelChannelIn_rData_rowEnd;
  wire                when_Stream_l368_2;
  wire                pixelChannelJoin_valid;
  wire                pixelChannelJoin_ready;
  wire       [7:0]    pixelChannelJoin_payload_0_pixel;
  wire                pixelChannelJoin_payload_0_frameStart;
  wire                pixelChannelJoin_payload_0_rowEnd;
  wire       [7:0]    pixelChannelJoin_payload_1_pixel;
  wire                pixelChannelJoin_payload_1_frameStart;
  wire                pixelChannelJoin_payload_1_rowEnd;
  wire       [7:0]    pixelChannelJoin_payload_2_pixel;
  wire                pixelChannelJoin_payload_2_frameStart;
  wire                pixelChannelJoin_payload_2_rowEnd;
  wire                pixelChannelJoin_fire;
  wire                pixelChannelJoin_fire_1;
  wire                pixelChannelJoin_fire_2;
  wire                pixelChannelJoin_translated_valid;
  wire                pixelChannelJoin_translated_ready;
  wire       [31:0]   pixelChannelJoin_translated_payload_pixel;
  wire                pixelChannelJoin_translated_payload_frameStart;
  wire                pixelChannelJoin_translated_payload_rowEnd;
  wire                pixelChannelJoin_translated_s2mPipe_valid;
  reg                 pixelChannelJoin_translated_s2mPipe_ready;
  wire       [31:0]   pixelChannelJoin_translated_s2mPipe_payload_pixel;
  wire                pixelChannelJoin_translated_s2mPipe_payload_frameStart;
  wire                pixelChannelJoin_translated_s2mPipe_payload_rowEnd;
  reg                 pixelChannelJoin_translated_rValid;
  reg        [31:0]   pixelChannelJoin_translated_rData_pixel;
  reg                 pixelChannelJoin_translated_rData_frameStart;
  reg                 pixelChannelJoin_translated_rData_rowEnd;
  wire                pixelChannelJoin_translated_s2mPipe_m2sPipe_valid;
  wire                pixelChannelJoin_translated_s2mPipe_m2sPipe_ready;
  wire       [31:0]   pixelChannelJoin_translated_s2mPipe_m2sPipe_payload_pixel;
  wire                pixelChannelJoin_translated_s2mPipe_m2sPipe_payload_frameStart;
  wire                pixelChannelJoin_translated_s2mPipe_m2sPipe_payload_rowEnd;
  reg                 pixelChannelJoin_translated_s2mPipe_rValid;
  reg        [31:0]   pixelChannelJoin_translated_s2mPipe_rData_pixel;
  reg                 pixelChannelJoin_translated_s2mPipe_rData_frameStart;
  reg                 pixelChannelJoin_translated_s2mPipe_rData_rowEnd;
  wire                when_Stream_l368_3;

  always @(*) begin
    bPixelChannelIn_ready = bPixelChannelIn_m2sPipe_ready;
    if(when_Stream_l368) begin
      bPixelChannelIn_ready = 1'b1;
    end
  end

  assign when_Stream_l368 = (! bPixelChannelIn_m2sPipe_valid);
  assign bPixelChannelIn_m2sPipe_valid = bPixelChannelIn_rValid;
  assign bPixelChannelIn_m2sPipe_payload_pixel = bPixelChannelIn_rData_pixel;
  assign bPixelChannelIn_m2sPipe_payload_frameStart = bPixelChannelIn_rData_frameStart;
  assign bPixelChannelIn_m2sPipe_payload_rowEnd = bPixelChannelIn_rData_rowEnd;
  always @(*) begin
    gPixelChannelIn_ready = gPixelChannelIn_m2sPipe_ready;
    if(when_Stream_l368_1) begin
      gPixelChannelIn_ready = 1'b1;
    end
  end

  assign when_Stream_l368_1 = (! gPixelChannelIn_m2sPipe_valid);
  assign gPixelChannelIn_m2sPipe_valid = gPixelChannelIn_rValid;
  assign gPixelChannelIn_m2sPipe_payload_pixel = gPixelChannelIn_rData_pixel;
  assign gPixelChannelIn_m2sPipe_payload_frameStart = gPixelChannelIn_rData_frameStart;
  assign gPixelChannelIn_m2sPipe_payload_rowEnd = gPixelChannelIn_rData_rowEnd;
  always @(*) begin
    rPixelChannelIn_ready = rPixelChannelIn_m2sPipe_ready;
    if(when_Stream_l368_2) begin
      rPixelChannelIn_ready = 1'b1;
    end
  end

  assign when_Stream_l368_2 = (! rPixelChannelIn_m2sPipe_valid);
  assign rPixelChannelIn_m2sPipe_valid = rPixelChannelIn_rValid;
  assign rPixelChannelIn_m2sPipe_payload_pixel = rPixelChannelIn_rData_pixel;
  assign rPixelChannelIn_m2sPipe_payload_frameStart = rPixelChannelIn_rData_frameStart;
  assign rPixelChannelIn_m2sPipe_payload_rowEnd = rPixelChannelIn_rData_rowEnd;
  assign pixelChannelJoin_payload_0_pixel = bPixelChannelIn_m2sPipe_payload_pixel;
  assign pixelChannelJoin_payload_0_frameStart = bPixelChannelIn_m2sPipe_payload_frameStart;
  assign pixelChannelJoin_payload_0_rowEnd = bPixelChannelIn_m2sPipe_payload_rowEnd;
  assign pixelChannelJoin_payload_1_pixel = gPixelChannelIn_m2sPipe_payload_pixel;
  assign pixelChannelJoin_payload_1_frameStart = gPixelChannelIn_m2sPipe_payload_frameStart;
  assign pixelChannelJoin_payload_1_rowEnd = gPixelChannelIn_m2sPipe_payload_rowEnd;
  assign pixelChannelJoin_payload_2_pixel = rPixelChannelIn_m2sPipe_payload_pixel;
  assign pixelChannelJoin_payload_2_frameStart = rPixelChannelIn_m2sPipe_payload_frameStart;
  assign pixelChannelJoin_payload_2_rowEnd = rPixelChannelIn_m2sPipe_payload_rowEnd;
  assign pixelChannelJoin_valid = ((bPixelChannelIn_m2sPipe_valid && gPixelChannelIn_m2sPipe_valid) && rPixelChannelIn_m2sPipe_valid);
  assign pixelChannelJoin_fire = (pixelChannelJoin_valid && pixelChannelJoin_ready);
  assign bPixelChannelIn_m2sPipe_ready = pixelChannelJoin_fire;
  assign pixelChannelJoin_fire_1 = (pixelChannelJoin_valid && pixelChannelJoin_ready);
  assign gPixelChannelIn_m2sPipe_ready = pixelChannelJoin_fire_1;
  assign pixelChannelJoin_fire_2 = (pixelChannelJoin_valid && pixelChannelJoin_ready);
  assign rPixelChannelIn_m2sPipe_ready = pixelChannelJoin_fire_2;
  assign pixelChannelJoin_translated_valid = pixelChannelJoin_valid;
  assign pixelChannelJoin_ready = pixelChannelJoin_translated_ready;
  assign pixelChannelJoin_translated_payload_pixel = {{{8'h0,pixelChannelJoin_payload_2_pixel},pixelChannelJoin_payload_1_pixel},pixelChannelJoin_payload_0_pixel};
  assign pixelChannelJoin_translated_payload_frameStart = pixelChannelJoin_payload_2_frameStart;
  assign pixelChannelJoin_translated_payload_rowEnd = pixelChannelJoin_payload_2_rowEnd;
  assign pixelChannelJoin_translated_ready = (! pixelChannelJoin_translated_rValid);
  assign pixelChannelJoin_translated_s2mPipe_valid = (pixelChannelJoin_translated_valid || pixelChannelJoin_translated_rValid);
  assign pixelChannelJoin_translated_s2mPipe_payload_pixel = (pixelChannelJoin_translated_rValid ? pixelChannelJoin_translated_rData_pixel : pixelChannelJoin_translated_payload_pixel);
  assign pixelChannelJoin_translated_s2mPipe_payload_frameStart = (pixelChannelJoin_translated_rValid ? pixelChannelJoin_translated_rData_frameStart : pixelChannelJoin_translated_payload_frameStart);
  assign pixelChannelJoin_translated_s2mPipe_payload_rowEnd = (pixelChannelJoin_translated_rValid ? pixelChannelJoin_translated_rData_rowEnd : pixelChannelJoin_translated_payload_rowEnd);
  always @(*) begin
    pixelChannelJoin_translated_s2mPipe_ready = pixelChannelJoin_translated_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_3) begin
      pixelChannelJoin_translated_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_3 = (! pixelChannelJoin_translated_s2mPipe_m2sPipe_valid);
  assign pixelChannelJoin_translated_s2mPipe_m2sPipe_valid = pixelChannelJoin_translated_s2mPipe_rValid;
  assign pixelChannelJoin_translated_s2mPipe_m2sPipe_payload_pixel = pixelChannelJoin_translated_s2mPipe_rData_pixel;
  assign pixelChannelJoin_translated_s2mPipe_m2sPipe_payload_frameStart = pixelChannelJoin_translated_s2mPipe_rData_frameStart;
  assign pixelChannelJoin_translated_s2mPipe_m2sPipe_payload_rowEnd = pixelChannelJoin_translated_s2mPipe_rData_rowEnd;
  assign allPixelChannelOut_valid = pixelChannelJoin_translated_s2mPipe_m2sPipe_valid;
  assign pixelChannelJoin_translated_s2mPipe_m2sPipe_ready = allPixelChannelOut_ready;
  assign allPixelChannelOut_payload_pixel = pixelChannelJoin_translated_s2mPipe_m2sPipe_payload_pixel;
  assign allPixelChannelOut_payload_frameStart = pixelChannelJoin_translated_s2mPipe_m2sPipe_payload_frameStart;
  assign allPixelChannelOut_payload_rowEnd = pixelChannelJoin_translated_s2mPipe_m2sPipe_payload_rowEnd;
  always @(posedge clk or negedge resetn) begin
    if(!resetn) begin
      bPixelChannelIn_rValid <= 1'b0;
      gPixelChannelIn_rValid <= 1'b0;
      rPixelChannelIn_rValid <= 1'b0;
      pixelChannelJoin_translated_rValid <= 1'b0;
      pixelChannelJoin_translated_s2mPipe_rValid <= 1'b0;
    end else begin
      if(bPixelChannelIn_ready) begin
        bPixelChannelIn_rValid <= bPixelChannelIn_valid;
      end
      if(gPixelChannelIn_ready) begin
        gPixelChannelIn_rValid <= gPixelChannelIn_valid;
      end
      if(rPixelChannelIn_ready) begin
        rPixelChannelIn_rValid <= rPixelChannelIn_valid;
      end
      if(pixelChannelJoin_translated_valid) begin
        pixelChannelJoin_translated_rValid <= 1'b1;
      end
      if(pixelChannelJoin_translated_s2mPipe_ready) begin
        pixelChannelJoin_translated_rValid <= 1'b0;
      end
      if(pixelChannelJoin_translated_s2mPipe_ready) begin
        pixelChannelJoin_translated_s2mPipe_rValid <= pixelChannelJoin_translated_s2mPipe_valid;
      end
    end
  end

  always @(posedge clk) begin
    if(bPixelChannelIn_ready) begin
      bPixelChannelIn_rData_pixel <= bPixelChannelIn_payload_pixel;
      bPixelChannelIn_rData_frameStart <= bPixelChannelIn_payload_frameStart;
      bPixelChannelIn_rData_rowEnd <= bPixelChannelIn_payload_rowEnd;
    end
    if(gPixelChannelIn_ready) begin
      gPixelChannelIn_rData_pixel <= gPixelChannelIn_payload_pixel;
      gPixelChannelIn_rData_frameStart <= gPixelChannelIn_payload_frameStart;
      gPixelChannelIn_rData_rowEnd <= gPixelChannelIn_payload_rowEnd;
    end
    if(rPixelChannelIn_ready) begin
      rPixelChannelIn_rData_pixel <= rPixelChannelIn_payload_pixel;
      rPixelChannelIn_rData_frameStart <= rPixelChannelIn_payload_frameStart;
      rPixelChannelIn_rData_rowEnd <= rPixelChannelIn_payload_rowEnd;
    end
    if(pixelChannelJoin_translated_ready) begin
      pixelChannelJoin_translated_rData_pixel <= pixelChannelJoin_translated_payload_pixel;
      pixelChannelJoin_translated_rData_frameStart <= pixelChannelJoin_translated_payload_frameStart;
      pixelChannelJoin_translated_rData_rowEnd <= pixelChannelJoin_translated_payload_rowEnd;
    end
    if(pixelChannelJoin_translated_s2mPipe_ready) begin
      pixelChannelJoin_translated_s2mPipe_rData_pixel <= pixelChannelJoin_translated_s2mPipe_payload_pixel;
      pixelChannelJoin_translated_s2mPipe_rData_frameStart <= pixelChannelJoin_translated_s2mPipe_payload_frameStart;
      pixelChannelJoin_translated_s2mPipe_rData_rowEnd <= pixelChannelJoin_translated_s2mPipe_payload_rowEnd;
    end
  end


endmodule

module SuperResolutionPart3_2 (
  input               pixelsIn_valid,
  output reg          pixelsIn_ready,
  input      [7:0]    pixelsIn_payload_pixel,
  input               pixelsIn_payload_frameStart,
  input               pixelsIn_payload_rowEnd,
  input               pixelsIn_payload_inpValid,
  input               startIn,
  output reg          pixelsOut_valid,
  input               pixelsOut_ready,
  output reg [7:0]    pixelsOut_payload_pixel,
  output reg          pixelsOut_payload_frameStart,
  output reg          pixelsOut_payload_rowEnd,
  output reg          inpThreeDoneOut,
  input      [7:0]    thresholdIn,
  input      [9:0]    widthIn,
  input      [9:0]    heightIn,
  input               clk,
  input               resetn
);
  localparam controlStateMachine_enumDef_8_BOOT = 2'd0;
  localparam controlStateMachine_enumDef_8_HOLD = 2'd1;
  localparam controlStateMachine_enumDef_8_PASS = 2'd2;
  localparam controlStateMachine_enumDef_8_EXTRA = 2'd3;

  reg        [7:0]    CICC1851_lineBufferOne_port1;
  reg        [7:0]    CICC1851_lineBufferOne_port2;
  reg        [7:0]    CICC1851_lineBufferTwo_port1;
  reg        [7:0]    CICC1851_lineBufferTwo_port2;
  reg        [7:0]    CICC1851_lineBufferThree_port1;
  reg        [7:0]    CICC1851_lineBufferThree_port2;
  reg        [0:0]    CICC1851_validBufferOne_port1;
  reg        [0:0]    CICC1851_validBufferOne_port2;
  reg        [0:0]    CICC1851_validBufferTwo_port1;
  reg        [0:0]    CICC1851_validBufferTwo_port2;
  reg        [0:0]    CICC1851_validBufferThree_port1;
  reg        [0:0]    CICC1851_validBufferThree_port2;
  wire                diffStage_controlPipe_fork_io_input_ready;
  wire                diffStage_controlPipe_fork_io_outputs_0_valid;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_frameStart;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_rowEnd;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_pipeValid;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_firstRow;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_lastRow;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_finalResult;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_mainCompare;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_counterCompare;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_horizontalCompare;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_verticalCompare;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_payload_mainDiff;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_payload_counterDiff;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_payload_horizontalDiff;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_payload_verticalDiff;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_isHorizontalMin;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_payload_minDiff;
  wire       [1:0]    diffStage_controlPipe_fork_io_outputs_0_payload_currentPosition;
  wire       [1:0]    diffStage_controlPipe_fork_io_outputs_0_payload_nextPosition;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_horizontalDirectionValid;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_verticalDirectionValid;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_mainDirectionValid;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_counterDirectionValid;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_inValidMinDiff;
  wire                diffStage_controlPipe_fork_io_outputs_1_valid;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_frameStart;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_rowEnd;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_pipeValid;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_firstRow;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_lastRow;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_finalResult;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_mainCompare;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_counterCompare;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_horizontalCompare;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_verticalCompare;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_1_payload_horizontalDiff;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_1_payload_verticalDiff;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_isHorizontalMin;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_1_payload_minDiff;
  wire       [1:0]    diffStage_controlPipe_fork_io_outputs_1_payload_currentPosition;
  wire       [1:0]    diffStage_controlPipe_fork_io_outputs_1_payload_nextPosition;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_horizontalDirectionValid;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_verticalDirectionValid;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_mainDirectionValid;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_counterDirectionValid;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_inValidMinDiff;
  wire       [11:0]   CICC1851_bufferRowCount_valueNext;
  wire       [0:0]    CICC1851_bufferRowCount_valueNext_1;
  wire       [11:0]   CICC1851_bufferWAddr_valueNext;
  wire       [0:0]    CICC1851_bufferWAddr_valueNext_1;
  wire       [11:0]   CICC1851_outPixelAddr_valueNext;
  wire       [0:0]    CICC1851_outPixelAddr_valueNext_1;
  wire       [11:0]   CICC1851_outRowCount_valueNext;
  wire       [0:0]    CICC1851_outRowCount_valueNext_1;
  wire       [11:0]   CICC1851_alreadySendRow_valueNext;
  wire       [0:0]    CICC1851_alreadySendRow_valueNext_1;
  wire       [11:0]   CICC1851_alreadySendCountInRow_valueNext;
  wire       [0:0]    CICC1851_alreadySendCountInRow_valueNext_1;
  wire       [0:0]    CICC1851_nextRowBuffer;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l226;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l226_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l226_2;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l227;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l227_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l227_2;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l270;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l270_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l270_2;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l271;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l271_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l271_2;
  wire       [7:0]    CICC1851_lineBufferOne_port;
  wire                CICC1851_lineBufferOne_port_1;
  wire       [7:0]    CICC1851_lineBufferTwo_port;
  wire                CICC1851_lineBufferTwo_port_1;
  wire       [7:0]    CICC1851_lineBufferThree_port;
  wire                CICC1851_lineBufferThree_port_1;
  wire       [0:0]    CICC1851_validBufferOne_port;
  wire                CICC1851_validBufferOne_port_1;
  wire       [0:0]    CICC1851_validBufferTwo_port;
  wire                CICC1851_validBufferTwo_port_1;
  wire       [0:0]    CICC1851_validBufferThree_port;
  wire                CICC1851_validBufferThree_port_1;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_1;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_2;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_3;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_4;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_5;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_6;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_7;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_8;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_9;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_10;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_11;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_12;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_13;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_14;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_15;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_16;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_17;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_18;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_19;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_20;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_21;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_22;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_23;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_24;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_25;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_26;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_27;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_28;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_29;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_30;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_31;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_32;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_33;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_34;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_35;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_36;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_37;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_38;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_39;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_40;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_41;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_42;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_43;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_44;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_45;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_46;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_47;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_48;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_49;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_50;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_51;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_52;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_53;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_54;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_55;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_56;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_57;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_58;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_59;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_60;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_61;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_62;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_63;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_64;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_65;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_66;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_67;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_68;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_69;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_70;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_71;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_72;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_73;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_74;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_75;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_76;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_77;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_78;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_79;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_80;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_81;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_82;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_83;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_84;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_85;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_86;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_87;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_88;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_89;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_90;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_91;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_92;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_93;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_94;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_95;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_96;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_97;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_98;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_99;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_100;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_101;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_102;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_103;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_104;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_105;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_106;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_107;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_108;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_109;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_110;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_111;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_112;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_113;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_114;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_115;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_116;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_117;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_118;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_119;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_120;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_121;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_122;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_123;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_124;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_125;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_126;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_127;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_128;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_129;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_130;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_131;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_132;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_133;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_134;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_135;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_136;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_137;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_138;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_139;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_140;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_141;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_142;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_143;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_144;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_145;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_146;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_147;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_148;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_149;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_150;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_151;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_152;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_153;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_154;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_155;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_156;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_157;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_158;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_159;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_160;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_161;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_162;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_163;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_164;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_165;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_166;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_167;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_168;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_169;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_170;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_171;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_172;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_173;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_174;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_175;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_176;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_177;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_178;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_179;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_180;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_181;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_182;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_183;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_184;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_185;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_186;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_187;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_188;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_189;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_190;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_191;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_192;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_193;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_194;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_195;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_196;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_197;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_198;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_199;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_200;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_201;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_202;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_203;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_204;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_205;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_206;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_207;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_208;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_209;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_210;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_211;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_212;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_213;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_214;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_215;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_216;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_217;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_218;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_219;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_220;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_221;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_222;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_223;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_224;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_225;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_226;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_227;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_228;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_229;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_230;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_231;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_232;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_233;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_234;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_235;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_236;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_237;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_238;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_239;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_240;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_241;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_242;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_243;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_244;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_245;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_246;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_247;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_248;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_249;
  wire       [11:0]   CICC1851_when_SuperResolutionPart3_l1202;
  wire       [11:0]   CICC1851_when_SuperResolutionPart3_l1205;
  wire       [11:0]   CICC1851_when_SuperResolutionPart3_l1205_1;
  wire       [11:0]   CICC1851_when_SuperResolutionPart3_l1205_2;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l1223;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l1223_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l1223_2;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l1224;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l1224_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l1224_2;
  reg                 inpThreeDone;
  reg                 startIn_regNext;
  wire                when_SuperResolutionPart3_l72;
  reg                 readDone;
  wire                when_SuperResolutionPart3_l75;
  reg                 startRead;
  wire                when_SuperResolutionPart3_l78;
  wire                when_SuperResolutionPart3_l78_1;
  reg                 frameStart;
  reg        [7:0]    inpThreshold;
  reg        [9:0]    bmpWidth;
  reg        [9:0]    bmpHeight;
  reg                 holdBuffer;
  wire                when_SuperResolutionPart3_l93;
  reg                 writeDone;
  wire                when_SuperResolutionPart3_l96;
  reg                 bufferRowCount_willIncrement;
  reg                 bufferRowCount_willClear;
  reg        [11:0]   bufferRowCount_valueNext;
  reg        [11:0]   bufferRowCount_value;
  wire                bufferRowCount_willOverflowIfInc;
  wire                bufferRowCount_willOverflow;
  reg                 bufferEnable;
  wire                when_SuperResolutionPart3_l102;
  wire                when_SuperResolutionPart3_l102_1;
  reg        [1:0]    bufferSwitch;
  reg        [1:0]    nextRowBuffer;
  reg        [1:0]    currentRowBuffer;
  reg                 bufferReuse;
  reg                 bufferWAddr_willIncrement;
  reg                 bufferWAddr_willClear;
  reg        [11:0]   bufferWAddr_valueNext;
  reg        [11:0]   bufferWAddr_value;
  wire                bufferWAddr_willOverflowIfInc;
  wire                bufferWAddr_willOverflow;
  reg                 outPixelAddr_willIncrement;
  reg                 outPixelAddr_willClear;
  reg        [11:0]   outPixelAddr_valueNext;
  reg        [11:0]   outPixelAddr_value;
  wire                outPixelAddr_willOverflowIfInc;
  wire                outPixelAddr_willOverflow;
  reg                 outRowCount_willIncrement;
  reg                 outRowCount_willClear;
  reg        [11:0]   outRowCount_valueNext;
  reg        [11:0]   outRowCount_value;
  wire                outRowCount_willOverflowIfInc;
  wire                outRowCount_willOverflow;
  reg                 alreadySendRow_willIncrement;
  reg                 alreadySendRow_willClear;
  reg        [11:0]   alreadySendRow_valueNext;
  reg        [11:0]   alreadySendRow_value;
  wire                alreadySendRow_willOverflowIfInc;
  wire                alreadySendRow_willOverflow;
  reg                 alreadySendCountInRow_willIncrement;
  reg                 alreadySendCountInRow_willClear;
  reg        [11:0]   alreadySendCountInRow_valueNext;
  reg        [11:0]   alreadySendCountInRow_value;
  wire                alreadySendCountInRow_willOverflowIfInc;
  wire                alreadySendCountInRow_willOverflow;
  reg                 alreadyReachRowEnd;
  reg                 alreadyReachFinalRow;
  reg                 outReachRowEnd;
  reg                 outReachFinalRow;
  reg                 bufferReachRowEnd;
  reg                 bufferReachFinalRow;
  reg        [7:0]    minDiff;
  reg        [7:0]    candidatePixel;
  reg                 isHorizontalDirection;
  reg                 inValidMinDiff;
  reg                 startIn_regNext_1;
  wire                when_SuperResolutionPart3_l154;
  reg        [11:0]   mainAddrOne;
  reg        [11:0]   counterAddrOne;
  reg        [11:0]   mainAddrTwo;
  reg        [11:0]   counterAddrTwo;
  reg        [11:0]   mainAddrThree;
  reg        [11:0]   counterAddrThree;
  wire                validStream_valid;
  reg                 validStream_ready;
  wire                controlStream_valid;
  wire                controlStream_ready;
  wire                controlStream_payload_frameStart;
  wire                controlStream_payload_rowEnd;
  wire                controlStream_payload_pipeValid;
  wire                controlStream_payload_firstRow;
  wire                controlStream_payload_lastRow;
  wire                controlStream_payload_finalResult;
  wire                controlStream_payload_mainCompare;
  wire                controlStream_payload_counterCompare;
  wire                controlStream_payload_horizontalCompare;
  wire                controlStream_payload_verticalCompare;
  wire       [7:0]    controlStream_payload_mainDiff;
  wire       [7:0]    controlStream_payload_counterDiff;
  wire       [7:0]    controlStream_payload_horizontalDiff;
  wire       [7:0]    controlStream_payload_verticalDiff;
  wire                controlStream_payload_isHorizontalMin;
  wire       [7:0]    controlStream_payload_minDiff;
  wire       [1:0]    controlStream_payload_currentPosition;
  wire       [1:0]    controlStream_payload_nextPosition;
  wire                controlStream_payload_horizontalDirectionValid;
  wire                controlStream_payload_verticalDirectionValid;
  wire                controlStream_payload_mainDirectionValid;
  wire                controlStream_payload_counterDirectionValid;
  wire                controlStream_payload_inValidMinDiff;
  reg                 controls_frameStart;
  reg                 controls_rowEnd;
  reg                 controls_pipeValid;
  reg                 controls_firstRow;
  reg                 controls_lastRow;
  reg                 controls_finalResult;
  wire                controls_mainCompare;
  wire                controls_counterCompare;
  wire                controls_horizontalCompare;
  wire                controls_verticalCompare;
  wire       [7:0]    controls_mainDiff;
  wire       [7:0]    controls_counterDiff;
  wire       [7:0]    controls_horizontalDiff;
  wire       [7:0]    controls_verticalDiff;
  wire                controls_isHorizontalMin;
  wire       [7:0]    controls_minDiff;
  reg        [1:0]    controls_currentPosition;
  reg        [1:0]    controls_nextPosition;
  wire                controls_horizontalDirectionValid;
  wire                controls_verticalDirectionValid;
  wire                controls_mainDirectionValid;
  wire                controls_counterDirectionValid;
  wire                controls_inValidMinDiff;
  wire       [59:0]   CICC1851_controls_frameStart;
  wire                mainPixelAddrOneStream_valid;
  wire                mainPixelAddrOneStream_ready;
  wire       [11:0]   mainPixelAddrOneStream_payload;
  wire                counterPixelAddrOneStream_valid;
  wire                counterPixelAddrOneStream_ready;
  wire       [11:0]   counterPixelAddrOneStream_payload;
  wire                mainPixelAddrTwoStream_valid;
  wire                mainPixelAddrTwoStream_ready;
  wire       [11:0]   mainPixelAddrTwoStream_payload;
  wire                counterPixelAddrTwoStream_valid;
  wire                counterPixelAddrTwoStream_ready;
  wire       [11:0]   counterPixelAddrTwoStream_payload;
  wire                mainPixelAddrThreeStream_valid;
  wire                mainPixelAddrThreeStream_ready;
  wire       [11:0]   mainPixelAddrThreeStream_payload;
  wire                counterPixelAddrThreeStream_valid;
  wire                counterPixelAddrThreeStream_ready;
  wire       [11:0]   counterPixelAddrThreeStream_payload;
  wire                mainValidAddrOneStream_valid;
  wire                mainValidAddrOneStream_ready;
  wire       [11:0]   mainValidAddrOneStream_payload;
  wire                counterValidAddrOneStream_valid;
  wire                counterValidAddrOneStream_ready;
  wire       [11:0]   counterValidAddrOneStream_payload;
  wire                mainValidAddrTwoStream_valid;
  wire                mainValidAddrTwoStream_ready;
  wire       [11:0]   mainValidAddrTwoStream_payload;
  wire                counterValidAddrTwoStream_valid;
  wire                counterValidAddrTwoStream_ready;
  wire       [11:0]   counterValidAddrTwoStream_payload;
  wire                mainValidAddrThreeStream_valid;
  wire                mainValidAddrThreeStream_ready;
  wire       [11:0]   mainValidAddrThreeStream_payload;
  wire                counterValidAddrThreeStream_valid;
  wire                counterValidAddrThreeStream_ready;
  wire       [11:0]   counterValidAddrThreeStream_payload;
  wire                pixelsIn_s2mPipe_valid;
  reg                 pixelsIn_s2mPipe_ready;
  wire       [7:0]    pixelsIn_s2mPipe_payload_pixel;
  wire                pixelsIn_s2mPipe_payload_frameStart;
  wire                pixelsIn_s2mPipe_payload_rowEnd;
  wire                pixelsIn_s2mPipe_payload_inpValid;
  reg                 pixelsIn_rValid;
  reg        [7:0]    pixelsIn_rData_pixel;
  reg                 pixelsIn_rData_frameStart;
  reg                 pixelsIn_rData_rowEnd;
  reg                 pixelsIn_rData_inpValid;
  wire                pixelsIn_s2mPipe_m2sPipe_valid;
  wire                pixelsIn_s2mPipe_m2sPipe_ready;
  wire       [7:0]    pixelsIn_s2mPipe_m2sPipe_payload_pixel;
  wire                pixelsIn_s2mPipe_m2sPipe_payload_frameStart;
  wire                pixelsIn_s2mPipe_m2sPipe_payload_rowEnd;
  wire                pixelsIn_s2mPipe_m2sPipe_payload_inpValid;
  reg                 pixelsIn_s2mPipe_rValid;
  reg        [7:0]    pixelsIn_s2mPipe_rData_pixel;
  reg                 pixelsIn_s2mPipe_rData_frameStart;
  reg                 pixelsIn_s2mPipe_rData_rowEnd;
  reg                 pixelsIn_s2mPipe_rData_inpValid;
  wire                when_Stream_l368;
  wire                passPixels_valid;
  wire                passPixels_ready;
  wire       [7:0]    passPixels_payload_pixel;
  wire                passPixels_payload_frameStart;
  wire                passPixels_payload_rowEnd;
  wire                passPixels_payload_inpValid;
  wire                passPixels_fire;
  wire                when_SuperResolutionPart3_l226;
  wire                passPixels_fire_1;
  wire                when_SuperResolutionPart3_l227;
  wire                passPixels_fire_2;
  wire                when_SuperResolutionPart3_l230;
  wire                passPixels_fire_3;
  wire                when_SuperResolutionPart3_l243;
  wire                when_SuperResolutionPart3_l244;
  wire                passPixels_fire_4;
  wire                when_SuperResolutionPart3_l251;
  wire                when_SuperResolutionPart3_l255;
  wire                passPixels_fire_5;
  wire                when_SuperResolutionPart3_l262;
  wire                pixelsOut_fire;
  wire                when_SuperResolutionPart3_l270;
  wire                pixelsOut_fire_1;
  wire                when_SuperResolutionPart3_l271;
  wire                pixelsOut_fire_2;
  wire                pixelsOut_fire_3;
  wire                when_SuperResolutionPart3_l282;
  wire                passPixels_fire_6;
  wire                passPixels_fire_7;
  wire                passPixels_fire_8;
  wire                passPixels_fire_9;
  wire                passPixels_fire_10;
  wire                passPixels_fire_11;
  wire                passPixels_fire_12;
  wire                mainPixelAddrOneStream_s2mPipe_valid;
  reg                 mainPixelAddrOneStream_s2mPipe_ready;
  wire       [11:0]   mainPixelAddrOneStream_s2mPipe_payload;
  reg                 mainPixelAddrOneStream_rValid;
  reg        [11:0]   mainPixelAddrOneStream_rData;
  wire                mainPixelAddrOneStream_s2mPipe_m2sPipe_valid;
  wire                mainPixelAddrOneStream_s2mPipe_m2sPipe_ready;
  wire       [11:0]   mainPixelAddrOneStream_s2mPipe_m2sPipe_payload;
  reg                 mainPixelAddrOneStream_s2mPipe_rValid;
  reg        [11:0]   mainPixelAddrOneStream_s2mPipe_rData;
  wire                when_Stream_l368_1;
  wire                CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_mainOnePixelStream_payload;
  reg                 CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_1;
  reg                 CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_mainOnePixelStream_payload_1;
  wire                readStage_mainOnePixelStream_valid;
  wire                readStage_mainOnePixelStream_ready;
  wire       [7:0]    readStage_mainOnePixelStream_payload;
  reg                 CICC1851_readStage_mainOnePixelStream_valid;
  reg        [7:0]    CICC1851_readStage_mainOnePixelStream_payload_2;
  wire                when_Stream_l368_2;
  wire                counterPixelAddrOneStream_s2mPipe_valid;
  reg                 counterPixelAddrOneStream_s2mPipe_ready;
  wire       [11:0]   counterPixelAddrOneStream_s2mPipe_payload;
  reg                 counterPixelAddrOneStream_rValid;
  reg        [11:0]   counterPixelAddrOneStream_rData;
  wire                counterPixelAddrOneStream_s2mPipe_m2sPipe_valid;
  wire                counterPixelAddrOneStream_s2mPipe_m2sPipe_ready;
  wire       [11:0]   counterPixelAddrOneStream_s2mPipe_m2sPipe_payload;
  reg                 counterPixelAddrOneStream_s2mPipe_rValid;
  reg        [11:0]   counterPixelAddrOneStream_s2mPipe_rData;
  wire                when_Stream_l368_3;
  wire                CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_counterOnePixelStream_payload;
  reg                 CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_2;
  reg                 CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_counterOnePixelStream_payload_1;
  wire                readStage_counterOnePixelStream_valid;
  wire                readStage_counterOnePixelStream_ready;
  wire       [7:0]    readStage_counterOnePixelStream_payload;
  reg                 CICC1851_readStage_counterOnePixelStream_valid;
  reg        [7:0]    CICC1851_readStage_counterOnePixelStream_payload_2;
  wire                when_Stream_l368_4;
  wire                mainPixelAddrTwoStream_s2mPipe_valid;
  reg                 mainPixelAddrTwoStream_s2mPipe_ready;
  wire       [11:0]   mainPixelAddrTwoStream_s2mPipe_payload;
  reg                 mainPixelAddrTwoStream_rValid;
  reg        [11:0]   mainPixelAddrTwoStream_rData;
  wire                mainPixelAddrTwoStream_s2mPipe_m2sPipe_valid;
  wire                mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire       [11:0]   mainPixelAddrTwoStream_s2mPipe_m2sPipe_payload;
  reg                 mainPixelAddrTwoStream_s2mPipe_rValid;
  reg        [11:0]   mainPixelAddrTwoStream_s2mPipe_rData;
  wire                when_Stream_l368_5;
  wire                CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_mainTwoPixelStream_payload;
  reg                 CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_3;
  reg                 CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_mainTwoPixelStream_payload_1;
  wire                readStage_mainTwoPixelStream_valid;
  wire                readStage_mainTwoPixelStream_ready;
  wire       [7:0]    readStage_mainTwoPixelStream_payload;
  reg                 CICC1851_readStage_mainTwoPixelStream_valid;
  reg        [7:0]    CICC1851_readStage_mainTwoPixelStream_payload_2;
  wire                when_Stream_l368_6;
  wire                counterPixelAddrTwoStream_s2mPipe_valid;
  reg                 counterPixelAddrTwoStream_s2mPipe_ready;
  wire       [11:0]   counterPixelAddrTwoStream_s2mPipe_payload;
  reg                 counterPixelAddrTwoStream_rValid;
  reg        [11:0]   counterPixelAddrTwoStream_rData;
  wire                counterPixelAddrTwoStream_s2mPipe_m2sPipe_valid;
  wire                counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire       [11:0]   counterPixelAddrTwoStream_s2mPipe_m2sPipe_payload;
  reg                 counterPixelAddrTwoStream_s2mPipe_rValid;
  reg        [11:0]   counterPixelAddrTwoStream_s2mPipe_rData;
  wire                when_Stream_l368_7;
  wire                CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_counterTwoPixelStream_payload;
  reg                 CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_4;
  reg                 CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_counterTwoPixelStream_payload_1;
  wire                readStage_counterTwoPixelStream_valid;
  wire                readStage_counterTwoPixelStream_ready;
  wire       [7:0]    readStage_counterTwoPixelStream_payload;
  reg                 CICC1851_readStage_counterTwoPixelStream_valid;
  reg        [7:0]    CICC1851_readStage_counterTwoPixelStream_payload_2;
  wire                when_Stream_l368_8;
  wire                mainPixelAddrThreeStream_s2mPipe_valid;
  reg                 mainPixelAddrThreeStream_s2mPipe_ready;
  wire       [11:0]   mainPixelAddrThreeStream_s2mPipe_payload;
  reg                 mainPixelAddrThreeStream_rValid;
  reg        [11:0]   mainPixelAddrThreeStream_rData;
  wire                mainPixelAddrThreeStream_s2mPipe_m2sPipe_valid;
  wire                mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready;
  wire       [11:0]   mainPixelAddrThreeStream_s2mPipe_m2sPipe_payload;
  reg                 mainPixelAddrThreeStream_s2mPipe_rValid;
  reg        [11:0]   mainPixelAddrThreeStream_s2mPipe_rData;
  wire                when_Stream_l368_9;
  wire                CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_mainThreePixelStream_payload;
  reg                 CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_5;
  reg                 CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_mainThreePixelStream_payload_1;
  wire                readStage_mainThreePixelStream_valid;
  wire                readStage_mainThreePixelStream_ready;
  wire       [7:0]    readStage_mainThreePixelStream_payload;
  reg                 CICC1851_readStage_mainThreePixelStream_valid;
  reg        [7:0]    CICC1851_readStage_mainThreePixelStream_payload_2;
  wire                when_Stream_l368_10;
  wire                counterPixelAddrThreeStream_s2mPipe_valid;
  reg                 counterPixelAddrThreeStream_s2mPipe_ready;
  wire       [11:0]   counterPixelAddrThreeStream_s2mPipe_payload;
  reg                 counterPixelAddrThreeStream_rValid;
  reg        [11:0]   counterPixelAddrThreeStream_rData;
  wire                counterPixelAddrThreeStream_s2mPipe_m2sPipe_valid;
  wire                counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready;
  wire       [11:0]   counterPixelAddrThreeStream_s2mPipe_m2sPipe_payload;
  reg                 counterPixelAddrThreeStream_s2mPipe_rValid;
  reg        [11:0]   counterPixelAddrThreeStream_s2mPipe_rData;
  wire                when_Stream_l368_11;
  wire                CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_counterThreePixelStream_payload;
  reg                 CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_6;
  reg                 CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_counterThreePixelStream_payload_1;
  wire                readStage_counterThreePixelStream_valid;
  wire                readStage_counterThreePixelStream_ready;
  wire       [7:0]    readStage_counterThreePixelStream_payload;
  reg                 CICC1851_readStage_counterThreePixelStream_valid;
  reg        [7:0]    CICC1851_readStage_counterThreePixelStream_payload_2;
  wire                when_Stream_l368_12;
  wire                mainValidAddrOneStream_s2mPipe_valid;
  reg                 mainValidAddrOneStream_s2mPipe_ready;
  wire       [11:0]   mainValidAddrOneStream_s2mPipe_payload;
  reg                 mainValidAddrOneStream_rValid;
  reg        [11:0]   mainValidAddrOneStream_rData;
  wire                mainValidAddrOneStream_s2mPipe_m2sPipe_valid;
  wire                mainValidAddrOneStream_s2mPipe_m2sPipe_ready;
  wire       [11:0]   mainValidAddrOneStream_s2mPipe_m2sPipe_payload;
  reg                 mainValidAddrOneStream_s2mPipe_rValid;
  reg        [11:0]   mainValidAddrOneStream_s2mPipe_rData;
  wire                when_Stream_l368_13;
  wire                CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_1;
  wire                CICC1851_readStage_mainOneValidStream_payload;
  reg                 CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_7;
  reg                 CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_3;
  reg                 CICC1851_readStage_mainOneValidStream_payload_1;
  wire                readStage_mainOneValidStream_valid;
  wire                readStage_mainOneValidStream_ready;
  wire                readStage_mainOneValidStream_payload;
  reg                 CICC1851_readStage_mainOneValidStream_valid;
  reg                 CICC1851_readStage_mainOneValidStream_payload_2;
  wire                when_Stream_l368_14;
  wire                counterValidAddrOneStream_s2mPipe_valid;
  reg                 counterValidAddrOneStream_s2mPipe_ready;
  wire       [11:0]   counterValidAddrOneStream_s2mPipe_payload;
  reg                 counterValidAddrOneStream_rValid;
  reg        [11:0]   counterValidAddrOneStream_rData;
  wire                counterValidAddrOneStream_s2mPipe_m2sPipe_valid;
  wire                counterValidAddrOneStream_s2mPipe_m2sPipe_ready;
  wire       [11:0]   counterValidAddrOneStream_s2mPipe_m2sPipe_payload;
  reg                 counterValidAddrOneStream_s2mPipe_rValid;
  reg        [11:0]   counterValidAddrOneStream_s2mPipe_rData;
  wire                when_Stream_l368_15;
  wire                CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_1;
  wire                CICC1851_readStage_counterOneValidStream_payload;
  reg                 CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_8;
  reg                 CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_3;
  reg                 CICC1851_readStage_counterOneValidStream_payload_1;
  wire                readStage_counterOneValidStream_valid;
  wire                readStage_counterOneValidStream_ready;
  wire                readStage_counterOneValidStream_payload;
  reg                 CICC1851_readStage_counterOneValidStream_valid;
  reg                 CICC1851_readStage_counterOneValidStream_payload_2;
  wire                when_Stream_l368_16;
  wire                mainValidAddrTwoStream_s2mPipe_valid;
  reg                 mainValidAddrTwoStream_s2mPipe_ready;
  wire       [11:0]   mainValidAddrTwoStream_s2mPipe_payload;
  reg                 mainValidAddrTwoStream_rValid;
  reg        [11:0]   mainValidAddrTwoStream_rData;
  wire                mainValidAddrTwoStream_s2mPipe_m2sPipe_valid;
  wire                mainValidAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire       [11:0]   mainValidAddrTwoStream_s2mPipe_m2sPipe_payload;
  reg                 mainValidAddrTwoStream_s2mPipe_rValid;
  reg        [11:0]   mainValidAddrTwoStream_s2mPipe_rData;
  wire                when_Stream_l368_17;
  wire                CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_1;
  wire                CICC1851_readStage_mainTwoValidStream_payload;
  reg                 CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_9;
  reg                 CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_3;
  reg                 CICC1851_readStage_mainTwoValidStream_payload_1;
  wire                readStage_mainTwoValidStream_valid;
  wire                readStage_mainTwoValidStream_ready;
  wire                readStage_mainTwoValidStream_payload;
  reg                 CICC1851_readStage_mainTwoValidStream_valid;
  reg                 CICC1851_readStage_mainTwoValidStream_payload_2;
  wire                when_Stream_l368_18;
  wire                counterValidAddrTwoStream_s2mPipe_valid;
  reg                 counterValidAddrTwoStream_s2mPipe_ready;
  wire       [11:0]   counterValidAddrTwoStream_s2mPipe_payload;
  reg                 counterValidAddrTwoStream_rValid;
  reg        [11:0]   counterValidAddrTwoStream_rData;
  wire                counterValidAddrTwoStream_s2mPipe_m2sPipe_valid;
  wire                counterValidAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire       [11:0]   counterValidAddrTwoStream_s2mPipe_m2sPipe_payload;
  reg                 counterValidAddrTwoStream_s2mPipe_rValid;
  reg        [11:0]   counterValidAddrTwoStream_s2mPipe_rData;
  wire                when_Stream_l368_19;
  wire                CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_1;
  wire                CICC1851_readStage_counterTwoValidStream_payload;
  reg                 CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_10;
  reg                 CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_3;
  reg                 CICC1851_readStage_counterTwoValidStream_payload_1;
  wire                readStage_counterTwoValidStream_valid;
  wire                readStage_counterTwoValidStream_ready;
  wire                readStage_counterTwoValidStream_payload;
  reg                 CICC1851_readStage_counterTwoValidStream_valid;
  reg                 CICC1851_readStage_counterTwoValidStream_payload_2;
  wire                when_Stream_l368_20;
  wire                mainValidAddrThreeStream_s2mPipe_valid;
  reg                 mainValidAddrThreeStream_s2mPipe_ready;
  wire       [11:0]   mainValidAddrThreeStream_s2mPipe_payload;
  reg                 mainValidAddrThreeStream_rValid;
  reg        [11:0]   mainValidAddrThreeStream_rData;
  wire                mainValidAddrThreeStream_s2mPipe_m2sPipe_valid;
  wire                mainValidAddrThreeStream_s2mPipe_m2sPipe_ready;
  wire       [11:0]   mainValidAddrThreeStream_s2mPipe_m2sPipe_payload;
  reg                 mainValidAddrThreeStream_s2mPipe_rValid;
  reg        [11:0]   mainValidAddrThreeStream_s2mPipe_rData;
  wire                when_Stream_l368_21;
  wire                CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_1;
  wire                CICC1851_readStage_mainThreeValidStream_payload;
  reg                 CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_11;
  reg                 CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_3;
  reg                 CICC1851_readStage_mainThreeValidStream_payload_1;
  wire                readStage_mainThreeValidStream_valid;
  wire                readStage_mainThreeValidStream_ready;
  wire                readStage_mainThreeValidStream_payload;
  reg                 CICC1851_readStage_mainThreeValidStream_valid;
  reg                 CICC1851_readStage_mainThreeValidStream_payload_2;
  wire                when_Stream_l368_22;
  wire                counterValidAddrThreeStream_s2mPipe_valid;
  reg                 counterValidAddrThreeStream_s2mPipe_ready;
  wire       [11:0]   counterValidAddrThreeStream_s2mPipe_payload;
  reg                 counterValidAddrThreeStream_rValid;
  reg        [11:0]   counterValidAddrThreeStream_rData;
  wire                counterValidAddrThreeStream_s2mPipe_m2sPipe_valid;
  wire                counterValidAddrThreeStream_s2mPipe_m2sPipe_ready;
  wire       [11:0]   counterValidAddrThreeStream_s2mPipe_m2sPipe_payload;
  reg                 counterValidAddrThreeStream_s2mPipe_rValid;
  reg        [11:0]   counterValidAddrThreeStream_s2mPipe_rData;
  wire                when_Stream_l368_23;
  wire                CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_1;
  wire                CICC1851_readStage_counterThreeValidStream_payload;
  reg                 CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_12;
  reg                 CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_3;
  reg                 CICC1851_readStage_counterThreeValidStream_payload_1;
  wire                readStage_counterThreeValidStream_valid;
  wire                readStage_counterThreeValidStream_ready;
  wire                readStage_counterThreeValidStream_payload;
  reg                 CICC1851_readStage_counterThreeValidStream_valid;
  reg                 CICC1851_readStage_counterThreeValidStream_payload_2;
  wire                when_Stream_l368_24;
  wire                controlStream_s2mPipe_valid;
  reg                 controlStream_s2mPipe_ready;
  wire                controlStream_s2mPipe_payload_frameStart;
  wire                controlStream_s2mPipe_payload_rowEnd;
  wire                controlStream_s2mPipe_payload_pipeValid;
  wire                controlStream_s2mPipe_payload_firstRow;
  wire                controlStream_s2mPipe_payload_lastRow;
  wire                controlStream_s2mPipe_payload_finalResult;
  wire                controlStream_s2mPipe_payload_mainCompare;
  wire                controlStream_s2mPipe_payload_counterCompare;
  wire                controlStream_s2mPipe_payload_horizontalCompare;
  wire                controlStream_s2mPipe_payload_verticalCompare;
  wire       [7:0]    controlStream_s2mPipe_payload_mainDiff;
  wire       [7:0]    controlStream_s2mPipe_payload_counterDiff;
  wire       [7:0]    controlStream_s2mPipe_payload_horizontalDiff;
  wire       [7:0]    controlStream_s2mPipe_payload_verticalDiff;
  wire                controlStream_s2mPipe_payload_isHorizontalMin;
  wire       [7:0]    controlStream_s2mPipe_payload_minDiff;
  wire       [1:0]    controlStream_s2mPipe_payload_currentPosition;
  wire       [1:0]    controlStream_s2mPipe_payload_nextPosition;
  wire                controlStream_s2mPipe_payload_horizontalDirectionValid;
  wire                controlStream_s2mPipe_payload_verticalDirectionValid;
  wire                controlStream_s2mPipe_payload_mainDirectionValid;
  wire                controlStream_s2mPipe_payload_counterDirectionValid;
  wire                controlStream_s2mPipe_payload_inValidMinDiff;
  reg                 controlStream_rValid;
  reg                 controlStream_rData_frameStart;
  reg                 controlStream_rData_rowEnd;
  reg                 controlStream_rData_pipeValid;
  reg                 controlStream_rData_firstRow;
  reg                 controlStream_rData_lastRow;
  reg                 controlStream_rData_finalResult;
  reg                 controlStream_rData_mainCompare;
  reg                 controlStream_rData_counterCompare;
  reg                 controlStream_rData_horizontalCompare;
  reg                 controlStream_rData_verticalCompare;
  reg        [7:0]    controlStream_rData_mainDiff;
  reg        [7:0]    controlStream_rData_counterDiff;
  reg        [7:0]    controlStream_rData_horizontalDiff;
  reg        [7:0]    controlStream_rData_verticalDiff;
  reg                 controlStream_rData_isHorizontalMin;
  reg        [7:0]    controlStream_rData_minDiff;
  reg        [1:0]    controlStream_rData_currentPosition;
  reg        [1:0]    controlStream_rData_nextPosition;
  reg                 controlStream_rData_horizontalDirectionValid;
  reg                 controlStream_rData_verticalDirectionValid;
  reg                 controlStream_rData_mainDirectionValid;
  reg                 controlStream_rData_counterDirectionValid;
  reg                 controlStream_rData_inValidMinDiff;
  wire                controlStream_s2mPipe_m2sPipe_valid;
  reg                 controlStream_s2mPipe_m2sPipe_ready;
  wire                controlStream_s2mPipe_m2sPipe_payload_frameStart;
  wire                controlStream_s2mPipe_m2sPipe_payload_rowEnd;
  wire                controlStream_s2mPipe_m2sPipe_payload_pipeValid;
  wire                controlStream_s2mPipe_m2sPipe_payload_firstRow;
  wire                controlStream_s2mPipe_m2sPipe_payload_lastRow;
  wire                controlStream_s2mPipe_m2sPipe_payload_finalResult;
  wire                controlStream_s2mPipe_m2sPipe_payload_mainCompare;
  wire                controlStream_s2mPipe_m2sPipe_payload_counterCompare;
  wire                controlStream_s2mPipe_m2sPipe_payload_horizontalCompare;
  wire                controlStream_s2mPipe_m2sPipe_payload_verticalCompare;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_payload_mainDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_payload_counterDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_payload_horizontalDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_payload_verticalDiff;
  wire                controlStream_s2mPipe_m2sPipe_payload_isHorizontalMin;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_payload_minDiff;
  wire       [1:0]    controlStream_s2mPipe_m2sPipe_payload_currentPosition;
  wire       [1:0]    controlStream_s2mPipe_m2sPipe_payload_nextPosition;
  wire                controlStream_s2mPipe_m2sPipe_payload_horizontalDirectionValid;
  wire                controlStream_s2mPipe_m2sPipe_payload_verticalDirectionValid;
  wire                controlStream_s2mPipe_m2sPipe_payload_mainDirectionValid;
  wire                controlStream_s2mPipe_m2sPipe_payload_counterDirectionValid;
  wire                controlStream_s2mPipe_m2sPipe_payload_inValidMinDiff;
  reg                 controlStream_s2mPipe_rValid;
  reg                 controlStream_s2mPipe_rData_frameStart;
  reg                 controlStream_s2mPipe_rData_rowEnd;
  reg                 controlStream_s2mPipe_rData_pipeValid;
  reg                 controlStream_s2mPipe_rData_firstRow;
  reg                 controlStream_s2mPipe_rData_lastRow;
  reg                 controlStream_s2mPipe_rData_finalResult;
  reg                 controlStream_s2mPipe_rData_mainCompare;
  reg                 controlStream_s2mPipe_rData_counterCompare;
  reg                 controlStream_s2mPipe_rData_horizontalCompare;
  reg                 controlStream_s2mPipe_rData_verticalCompare;
  reg        [7:0]    controlStream_s2mPipe_rData_mainDiff;
  reg        [7:0]    controlStream_s2mPipe_rData_counterDiff;
  reg        [7:0]    controlStream_s2mPipe_rData_horizontalDiff;
  reg        [7:0]    controlStream_s2mPipe_rData_verticalDiff;
  reg                 controlStream_s2mPipe_rData_isHorizontalMin;
  reg        [7:0]    controlStream_s2mPipe_rData_minDiff;
  reg        [1:0]    controlStream_s2mPipe_rData_currentPosition;
  reg        [1:0]    controlStream_s2mPipe_rData_nextPosition;
  reg                 controlStream_s2mPipe_rData_horizontalDirectionValid;
  reg                 controlStream_s2mPipe_rData_verticalDirectionValid;
  reg                 controlStream_s2mPipe_rData_mainDirectionValid;
  reg                 controlStream_s2mPipe_rData_counterDirectionValid;
  reg                 controlStream_s2mPipe_rData_inValidMinDiff;
  wire                when_Stream_l368_25;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_valid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_ready;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_frameStart;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_rowEnd;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_pipeValid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_firstRow;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_lastRow;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_finalResult;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainCompare;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterCompare;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_horizontalCompare;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_verticalCompare;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_horizontalDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_verticalDiff;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_isHorizontalMin;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_minDiff;
  wire       [1:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_currentPosition;
  wire       [1:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_nextPosition;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_horizontalDirectionValid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_verticalDirectionValid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDirectionValid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDirectionValid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_inValidMinDiff;
  reg                 controlStream_s2mPipe_m2sPipe_rValid;
  reg                 controlStream_s2mPipe_m2sPipe_rData_frameStart;
  reg                 controlStream_s2mPipe_m2sPipe_rData_rowEnd;
  reg                 controlStream_s2mPipe_m2sPipe_rData_pipeValid;
  reg                 controlStream_s2mPipe_m2sPipe_rData_firstRow;
  reg                 controlStream_s2mPipe_m2sPipe_rData_lastRow;
  reg                 controlStream_s2mPipe_m2sPipe_rData_finalResult;
  reg                 controlStream_s2mPipe_m2sPipe_rData_mainCompare;
  reg                 controlStream_s2mPipe_m2sPipe_rData_counterCompare;
  reg                 controlStream_s2mPipe_m2sPipe_rData_horizontalCompare;
  reg                 controlStream_s2mPipe_m2sPipe_rData_verticalCompare;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_rData_mainDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_rData_counterDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_rData_horizontalDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_rData_verticalDiff;
  reg                 controlStream_s2mPipe_m2sPipe_rData_isHorizontalMin;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_rData_minDiff;
  reg        [1:0]    controlStream_s2mPipe_m2sPipe_rData_currentPosition;
  reg        [1:0]    controlStream_s2mPipe_m2sPipe_rData_nextPosition;
  reg                 controlStream_s2mPipe_m2sPipe_rData_horizontalDirectionValid;
  reg                 controlStream_s2mPipe_m2sPipe_rData_verticalDirectionValid;
  reg                 controlStream_s2mPipe_m2sPipe_rData_mainDirectionValid;
  reg                 controlStream_s2mPipe_m2sPipe_rData_counterDirectionValid;
  reg                 controlStream_s2mPipe_m2sPipe_rData_inValidMinDiff;
  wire                when_Stream_l368_26;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_valid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_frameStart;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_rowEnd;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_pipeValid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_firstRow;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_lastRow;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_finalResult;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainCompare;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterCompare;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_horizontalCompare;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_verticalCompare;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_horizontalDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_verticalDiff;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_isHorizontalMin;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_minDiff;
  wire       [1:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_currentPosition;
  wire       [1:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_nextPosition;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_horizontalDirectionValid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_verticalDirectionValid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainDirectionValid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterDirectionValid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_inValidMinDiff;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_frameStart;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_rowEnd;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_pipeValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_firstRow;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_lastRow;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_finalResult;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainCompare;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterCompare;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_horizontalCompare;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_verticalCompare;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_horizontalDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_verticalDiff;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_isHorizontalMin;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_minDiff;
  reg        [1:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_currentPosition;
  reg        [1:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_nextPosition;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_horizontalDirectionValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_verticalDirectionValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainDirectionValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterDirectionValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_inValidMinDiff;
  wire                readStage_controlPipe_valid;
  wire                readStage_controlPipe_ready;
  wire                readStage_controlPipe_payload_frameStart;
  wire                readStage_controlPipe_payload_rowEnd;
  wire                readStage_controlPipe_payload_pipeValid;
  wire                readStage_controlPipe_payload_firstRow;
  wire                readStage_controlPipe_payload_lastRow;
  wire                readStage_controlPipe_payload_finalResult;
  wire                readStage_controlPipe_payload_mainCompare;
  wire                readStage_controlPipe_payload_counterCompare;
  wire                readStage_controlPipe_payload_horizontalCompare;
  wire                readStage_controlPipe_payload_verticalCompare;
  wire       [7:0]    readStage_controlPipe_payload_mainDiff;
  wire       [7:0]    readStage_controlPipe_payload_counterDiff;
  wire       [7:0]    readStage_controlPipe_payload_horizontalDiff;
  wire       [7:0]    readStage_controlPipe_payload_verticalDiff;
  wire                readStage_controlPipe_payload_isHorizontalMin;
  wire       [7:0]    readStage_controlPipe_payload_minDiff;
  wire       [1:0]    readStage_controlPipe_payload_currentPosition;
  wire       [1:0]    readStage_controlPipe_payload_nextPosition;
  wire                readStage_controlPipe_payload_horizontalDirectionValid;
  wire                readStage_controlPipe_payload_verticalDirectionValid;
  wire                readStage_controlPipe_payload_mainDirectionValid;
  wire                readStage_controlPipe_payload_counterDirectionValid;
  wire                readStage_controlPipe_payload_inValidMinDiff;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_frameStart;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_rowEnd;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_pipeValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_firstRow;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_lastRow;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_finalResult;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainCompare;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterCompare;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_horizontalCompare;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_verticalCompare;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_horizontalDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_verticalDiff;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_isHorizontalMin;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_minDiff;
  reg        [1:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_currentPosition;
  reg        [1:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_nextPosition;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_horizontalDirectionValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_verticalDirectionValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainDirectionValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterDirectionValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_inValidMinDiff;
  wire                when_Stream_l368_27;
  wire                readStage_mainOnePixelStream_s2mPipe_valid;
  reg                 readStage_mainOnePixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_mainOnePixelStream_s2mPipe_payload;
  reg                 readStage_mainOnePixelStream_rValid;
  reg        [7:0]    readStage_mainOnePixelStream_rData;
  wire                compareStage_mainOnePixelStream_valid;
  wire                compareStage_mainOnePixelStream_ready;
  wire       [7:0]    compareStage_mainOnePixelStream_payload;
  reg                 readStage_mainOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_mainOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_28;
  wire                readStage_counterOnePixelStream_s2mPipe_valid;
  reg                 readStage_counterOnePixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_counterOnePixelStream_s2mPipe_payload;
  reg                 readStage_counterOnePixelStream_rValid;
  reg        [7:0]    readStage_counterOnePixelStream_rData;
  wire                compareStage_counterOnePixelStream_valid;
  wire                compareStage_counterOnePixelStream_ready;
  wire       [7:0]    compareStage_counterOnePixelStream_payload;
  reg                 readStage_counterOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_counterOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_29;
  wire                readStage_mainTwoPixelStream_s2mPipe_valid;
  reg                 readStage_mainTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_mainTwoPixelStream_s2mPipe_payload;
  reg                 readStage_mainTwoPixelStream_rValid;
  reg        [7:0]    readStage_mainTwoPixelStream_rData;
  wire                compareStage_mainTwoPixelStream_valid;
  wire                compareStage_mainTwoPixelStream_ready;
  wire       [7:0]    compareStage_mainTwoPixelStream_payload;
  reg                 readStage_mainTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_mainTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_30;
  wire                readStage_counterTwoPixelStream_s2mPipe_valid;
  reg                 readStage_counterTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_counterTwoPixelStream_s2mPipe_payload;
  reg                 readStage_counterTwoPixelStream_rValid;
  reg        [7:0]    readStage_counterTwoPixelStream_rData;
  wire                compareStage_counterTwoPixelStream_valid;
  wire                compareStage_counterTwoPixelStream_ready;
  wire       [7:0]    compareStage_counterTwoPixelStream_payload;
  reg                 readStage_counterTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_counterTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_31;
  wire                readStage_mainThreePixelStream_s2mPipe_valid;
  reg                 readStage_mainThreePixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_mainThreePixelStream_s2mPipe_payload;
  reg                 readStage_mainThreePixelStream_rValid;
  reg        [7:0]    readStage_mainThreePixelStream_rData;
  wire                compareStage_mainThreePixelStream_valid;
  wire                compareStage_mainThreePixelStream_ready;
  wire       [7:0]    compareStage_mainThreePixelStream_payload;
  reg                 readStage_mainThreePixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_mainThreePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_32;
  wire                readStage_counterThreePixelStream_s2mPipe_valid;
  reg                 readStage_counterThreePixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_counterThreePixelStream_s2mPipe_payload;
  reg                 readStage_counterThreePixelStream_rValid;
  reg        [7:0]    readStage_counterThreePixelStream_rData;
  wire                compareStage_counterThreePixelStream_valid;
  wire                compareStage_counterThreePixelStream_ready;
  wire       [7:0]    compareStage_counterThreePixelStream_payload;
  reg                 readStage_counterThreePixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_counterThreePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_33;
  wire                readStage_mainOneValidStream_s2mPipe_valid;
  reg                 readStage_mainOneValidStream_s2mPipe_ready;
  wire                readStage_mainOneValidStream_s2mPipe_payload;
  reg                 readStage_mainOneValidStream_rValid;
  reg                 readStage_mainOneValidStream_rData;
  wire                compareStage_mainOneValidStream_valid;
  wire                compareStage_mainOneValidStream_ready;
  wire                compareStage_mainOneValidStream_payload;
  reg                 readStage_mainOneValidStream_s2mPipe_rValid;
  reg                 readStage_mainOneValidStream_s2mPipe_rData;
  wire                when_Stream_l368_34;
  wire                readStage_counterOneValidStream_s2mPipe_valid;
  reg                 readStage_counterOneValidStream_s2mPipe_ready;
  wire                readStage_counterOneValidStream_s2mPipe_payload;
  reg                 readStage_counterOneValidStream_rValid;
  reg                 readStage_counterOneValidStream_rData;
  wire                compareStage_counterOneValidStream_valid;
  wire                compareStage_counterOneValidStream_ready;
  wire                compareStage_counterOneValidStream_payload;
  reg                 readStage_counterOneValidStream_s2mPipe_rValid;
  reg                 readStage_counterOneValidStream_s2mPipe_rData;
  wire                when_Stream_l368_35;
  wire                readStage_mainTwoValidStream_s2mPipe_valid;
  reg                 readStage_mainTwoValidStream_s2mPipe_ready;
  wire                readStage_mainTwoValidStream_s2mPipe_payload;
  reg                 readStage_mainTwoValidStream_rValid;
  reg                 readStage_mainTwoValidStream_rData;
  wire                compareStage_mainTwoValidStream_valid;
  wire                compareStage_mainTwoValidStream_ready;
  wire                compareStage_mainTwoValidStream_payload;
  reg                 readStage_mainTwoValidStream_s2mPipe_rValid;
  reg                 readStage_mainTwoValidStream_s2mPipe_rData;
  wire                when_Stream_l368_36;
  wire                readStage_counterTwoValidStream_s2mPipe_valid;
  reg                 readStage_counterTwoValidStream_s2mPipe_ready;
  wire                readStage_counterTwoValidStream_s2mPipe_payload;
  reg                 readStage_counterTwoValidStream_rValid;
  reg                 readStage_counterTwoValidStream_rData;
  wire                compareStage_counterTwoValidStream_valid;
  wire                compareStage_counterTwoValidStream_ready;
  wire                compareStage_counterTwoValidStream_payload;
  reg                 readStage_counterTwoValidStream_s2mPipe_rValid;
  reg                 readStage_counterTwoValidStream_s2mPipe_rData;
  wire                when_Stream_l368_37;
  wire                readStage_mainThreeValidStream_s2mPipe_valid;
  reg                 readStage_mainThreeValidStream_s2mPipe_ready;
  wire                readStage_mainThreeValidStream_s2mPipe_payload;
  reg                 readStage_mainThreeValidStream_rValid;
  reg                 readStage_mainThreeValidStream_rData;
  wire                compareStage_mainThreeValidStream_valid;
  wire                compareStage_mainThreeValidStream_ready;
  wire                compareStage_mainThreeValidStream_payload;
  reg                 readStage_mainThreeValidStream_s2mPipe_rValid;
  reg                 readStage_mainThreeValidStream_s2mPipe_rData;
  wire                when_Stream_l368_38;
  wire                readStage_counterThreeValidStream_s2mPipe_valid;
  reg                 readStage_counterThreeValidStream_s2mPipe_ready;
  wire                readStage_counterThreeValidStream_s2mPipe_payload;
  reg                 readStage_counterThreeValidStream_rValid;
  reg                 readStage_counterThreeValidStream_rData;
  wire                compareStage_counterThreeValidStream_valid;
  wire                compareStage_counterThreeValidStream_ready;
  wire                compareStage_counterThreeValidStream_payload;
  reg                 readStage_counterThreeValidStream_s2mPipe_rValid;
  reg                 readStage_counterThreeValidStream_s2mPipe_rData;
  wire                when_Stream_l368_39;
  reg                 CICC1851_readStage_controlPipe_translated_payload_mainCompare;
  reg                 CICC1851_readStage_controlPipe_translated_payload_counterCompare;
  reg                 CICC1851_readStage_controlPipe_translated_payload_horizontalCompare;
  reg                 CICC1851_readStage_controlPipe_translated_payload_verticalCompare;
  reg                 CICC1851_readStage_controlPipe_translated_payload_horizontalDirectionValid;
  reg                 CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid;
  reg                 CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid;
  reg                 CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid;
  wire                when_SuperResolutionPart3_l342;
  wire                when_SuperResolutionPart3_l344;
  wire                when_SuperResolutionPart3_l345;
  wire                when_SuperResolutionPart3_l348;
  wire                when_SuperResolutionPart3_l351;
  wire                when_SuperResolutionPart3_l347;
  wire                when_SuperResolutionPart3_l356;
  wire                when_SuperResolutionPart3_l357;
  wire                when_SuperResolutionPart3_l365;
  wire                when_SuperResolutionPart3_l373;
  wire                when_SuperResolutionPart3_l378;
  wire                when_SuperResolutionPart3_l383;
  wire                when_SuperResolutionPart3_l391;
  wire                when_SuperResolutionPart3_l396;
  wire                when_SuperResolutionPart3_l401;
  wire                when_SuperResolutionPart3_l409;
  wire                when_SuperResolutionPart3_l377;
  wire                when_SuperResolutionPart3_l415;
  wire                when_SuperResolutionPart3_l416;
  wire                when_SuperResolutionPart3_l419;
  wire                when_SuperResolutionPart3_l422;
  wire                when_SuperResolutionPart3_l424;
  wire                when_SuperResolutionPart3_l432;
  wire                when_SuperResolutionPart3_l441;
  wire                when_SuperResolutionPart3_l449;
  wire                when_SuperResolutionPart3_l458;
  wire                when_SuperResolutionPart3_l460;
  wire                when_SuperResolutionPart3_l463;
  wire                when_SuperResolutionPart3_l465;
  wire                when_SuperResolutionPart3_l470;
  wire                when_SuperResolutionPart3_l477;
  wire                when_SuperResolutionPart3_l485;
  wire                when_SuperResolutionPart3_l487;
  wire                when_SuperResolutionPart3_l490;
  wire                when_SuperResolutionPart3_l492;
  wire                when_SuperResolutionPart3_l497;
  wire                when_SuperResolutionPart3_l500;
  wire                when_SuperResolutionPart3_l502;
  wire                when_SuperResolutionPart3_l504;
  wire                when_SuperResolutionPart3_l511;
  wire                when_SuperResolutionPart3_l519;
  wire                when_SuperResolutionPart3_l521;
  wire                when_SuperResolutionPart3_l524;
  wire                when_SuperResolutionPart3_l526;
  wire                when_SuperResolutionPart3_l531;
  wire                when_SuperResolutionPart3_l539;
  wire                when_SuperResolutionPart3_l547;
  wire                when_SuperResolutionPart3_l549;
  wire                when_SuperResolutionPart3_l552;
  wire                when_SuperResolutionPart3_l554;
  wire                when_SuperResolutionPart3_l559;
  wire                when_SuperResolutionPart3_l562;
  wire                when_SuperResolutionPart3_l564;
  wire                when_SuperResolutionPart3_l566;
  wire                when_SuperResolutionPart3_l573;
  wire                when_SuperResolutionPart3_l581;
  wire                when_SuperResolutionPart3_l583;
  wire                when_SuperResolutionPart3_l586;
  wire                when_SuperResolutionPart3_l588;
  wire                when_SuperResolutionPart3_l593;
  wire                when_SuperResolutionPart3_l601;
  wire                when_SuperResolutionPart3_l609;
  wire                when_SuperResolutionPart3_l611;
  wire                when_SuperResolutionPart3_l614;
  wire                when_SuperResolutionPart3_l616;
  wire                when_SuperResolutionPart3_l496;
  wire                readStage_controlPipe_translated_valid;
  wire                readStage_controlPipe_translated_ready;
  wire                readStage_controlPipe_translated_payload_frameStart;
  wire                readStage_controlPipe_translated_payload_rowEnd;
  wire                readStage_controlPipe_translated_payload_pipeValid;
  wire                readStage_controlPipe_translated_payload_firstRow;
  wire                readStage_controlPipe_translated_payload_lastRow;
  wire                readStage_controlPipe_translated_payload_finalResult;
  wire                readStage_controlPipe_translated_payload_mainCompare;
  wire                readStage_controlPipe_translated_payload_counterCompare;
  wire                readStage_controlPipe_translated_payload_horizontalCompare;
  wire                readStage_controlPipe_translated_payload_verticalCompare;
  wire       [7:0]    readStage_controlPipe_translated_payload_mainDiff;
  wire       [7:0]    readStage_controlPipe_translated_payload_counterDiff;
  wire       [7:0]    readStage_controlPipe_translated_payload_horizontalDiff;
  wire       [7:0]    readStage_controlPipe_translated_payload_verticalDiff;
  wire                readStage_controlPipe_translated_payload_isHorizontalMin;
  wire       [7:0]    readStage_controlPipe_translated_payload_minDiff;
  wire       [1:0]    readStage_controlPipe_translated_payload_currentPosition;
  wire       [1:0]    readStage_controlPipe_translated_payload_nextPosition;
  wire                readStage_controlPipe_translated_payload_horizontalDirectionValid;
  wire                readStage_controlPipe_translated_payload_verticalDirectionValid;
  wire                readStage_controlPipe_translated_payload_mainDirectionValid;
  wire                readStage_controlPipe_translated_payload_counterDirectionValid;
  wire                readStage_controlPipe_translated_payload_inValidMinDiff;
  wire                readStage_controlPipe_translated_s2mPipe_valid;
  reg                 readStage_controlPipe_translated_s2mPipe_ready;
  wire                readStage_controlPipe_translated_s2mPipe_payload_frameStart;
  wire                readStage_controlPipe_translated_s2mPipe_payload_rowEnd;
  wire                readStage_controlPipe_translated_s2mPipe_payload_pipeValid;
  wire                readStage_controlPipe_translated_s2mPipe_payload_firstRow;
  wire                readStage_controlPipe_translated_s2mPipe_payload_lastRow;
  wire                readStage_controlPipe_translated_s2mPipe_payload_finalResult;
  wire                readStage_controlPipe_translated_s2mPipe_payload_mainCompare;
  wire                readStage_controlPipe_translated_s2mPipe_payload_counterCompare;
  wire                readStage_controlPipe_translated_s2mPipe_payload_horizontalCompare;
  wire                readStage_controlPipe_translated_s2mPipe_payload_verticalCompare;
  wire       [7:0]    readStage_controlPipe_translated_s2mPipe_payload_mainDiff;
  wire       [7:0]    readStage_controlPipe_translated_s2mPipe_payload_counterDiff;
  wire       [7:0]    readStage_controlPipe_translated_s2mPipe_payload_horizontalDiff;
  wire       [7:0]    readStage_controlPipe_translated_s2mPipe_payload_verticalDiff;
  wire                readStage_controlPipe_translated_s2mPipe_payload_isHorizontalMin;
  wire       [7:0]    readStage_controlPipe_translated_s2mPipe_payload_minDiff;
  wire       [1:0]    readStage_controlPipe_translated_s2mPipe_payload_currentPosition;
  wire       [1:0]    readStage_controlPipe_translated_s2mPipe_payload_nextPosition;
  wire                readStage_controlPipe_translated_s2mPipe_payload_horizontalDirectionValid;
  wire                readStage_controlPipe_translated_s2mPipe_payload_verticalDirectionValid;
  wire                readStage_controlPipe_translated_s2mPipe_payload_mainDirectionValid;
  wire                readStage_controlPipe_translated_s2mPipe_payload_counterDirectionValid;
  wire                readStage_controlPipe_translated_s2mPipe_payload_inValidMinDiff;
  reg                 readStage_controlPipe_translated_rValid;
  reg                 readStage_controlPipe_translated_rData_frameStart;
  reg                 readStage_controlPipe_translated_rData_rowEnd;
  reg                 readStage_controlPipe_translated_rData_pipeValid;
  reg                 readStage_controlPipe_translated_rData_firstRow;
  reg                 readStage_controlPipe_translated_rData_lastRow;
  reg                 readStage_controlPipe_translated_rData_finalResult;
  reg                 readStage_controlPipe_translated_rData_mainCompare;
  reg                 readStage_controlPipe_translated_rData_counterCompare;
  reg                 readStage_controlPipe_translated_rData_horizontalCompare;
  reg                 readStage_controlPipe_translated_rData_verticalCompare;
  reg        [7:0]    readStage_controlPipe_translated_rData_mainDiff;
  reg        [7:0]    readStage_controlPipe_translated_rData_counterDiff;
  reg        [7:0]    readStage_controlPipe_translated_rData_horizontalDiff;
  reg        [7:0]    readStage_controlPipe_translated_rData_verticalDiff;
  reg                 readStage_controlPipe_translated_rData_isHorizontalMin;
  reg        [7:0]    readStage_controlPipe_translated_rData_minDiff;
  reg        [1:0]    readStage_controlPipe_translated_rData_currentPosition;
  reg        [1:0]    readStage_controlPipe_translated_rData_nextPosition;
  reg                 readStage_controlPipe_translated_rData_horizontalDirectionValid;
  reg                 readStage_controlPipe_translated_rData_verticalDirectionValid;
  reg                 readStage_controlPipe_translated_rData_mainDirectionValid;
  reg                 readStage_controlPipe_translated_rData_counterDirectionValid;
  reg                 readStage_controlPipe_translated_rData_inValidMinDiff;
  wire                compareStage_controlPipe_valid;
  wire                compareStage_controlPipe_ready;
  wire                compareStage_controlPipe_payload_frameStart;
  wire                compareStage_controlPipe_payload_rowEnd;
  wire                compareStage_controlPipe_payload_pipeValid;
  wire                compareStage_controlPipe_payload_firstRow;
  wire                compareStage_controlPipe_payload_lastRow;
  wire                compareStage_controlPipe_payload_finalResult;
  wire                compareStage_controlPipe_payload_mainCompare;
  wire                compareStage_controlPipe_payload_counterCompare;
  wire                compareStage_controlPipe_payload_horizontalCompare;
  wire                compareStage_controlPipe_payload_verticalCompare;
  wire       [7:0]    compareStage_controlPipe_payload_mainDiff;
  wire       [7:0]    compareStage_controlPipe_payload_counterDiff;
  wire       [7:0]    compareStage_controlPipe_payload_horizontalDiff;
  wire       [7:0]    compareStage_controlPipe_payload_verticalDiff;
  wire                compareStage_controlPipe_payload_isHorizontalMin;
  wire       [7:0]    compareStage_controlPipe_payload_minDiff;
  wire       [1:0]    compareStage_controlPipe_payload_currentPosition;
  wire       [1:0]    compareStage_controlPipe_payload_nextPosition;
  wire                compareStage_controlPipe_payload_horizontalDirectionValid;
  wire                compareStage_controlPipe_payload_verticalDirectionValid;
  wire                compareStage_controlPipe_payload_mainDirectionValid;
  wire                compareStage_controlPipe_payload_counterDirectionValid;
  wire                compareStage_controlPipe_payload_inValidMinDiff;
  reg                 readStage_controlPipe_translated_s2mPipe_rValid;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_frameStart;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_rowEnd;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_pipeValid;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_firstRow;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_lastRow;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_finalResult;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_mainCompare;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_counterCompare;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_horizontalCompare;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_verticalCompare;
  reg        [7:0]    readStage_controlPipe_translated_s2mPipe_rData_mainDiff;
  reg        [7:0]    readStage_controlPipe_translated_s2mPipe_rData_counterDiff;
  reg        [7:0]    readStage_controlPipe_translated_s2mPipe_rData_horizontalDiff;
  reg        [7:0]    readStage_controlPipe_translated_s2mPipe_rData_verticalDiff;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_isHorizontalMin;
  reg        [7:0]    readStage_controlPipe_translated_s2mPipe_rData_minDiff;
  reg        [1:0]    readStage_controlPipe_translated_s2mPipe_rData_currentPosition;
  reg        [1:0]    readStage_controlPipe_translated_s2mPipe_rData_nextPosition;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_horizontalDirectionValid;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_verticalDirectionValid;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_mainDirectionValid;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_counterDirectionValid;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_inValidMinDiff;
  wire                when_Stream_l368_40;
  wire                compareStage_mainOnePixelStream_s2mPipe_valid;
  reg                 compareStage_mainOnePixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_mainOnePixelStream_s2mPipe_payload;
  reg                 compareStage_mainOnePixelStream_rValid;
  reg        [7:0]    compareStage_mainOnePixelStream_rData;
  wire                diffStage_mainOnePixelStream_valid;
  wire                diffStage_mainOnePixelStream_ready;
  wire       [7:0]    diffStage_mainOnePixelStream_payload;
  reg                 compareStage_mainOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_mainOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_41;
  wire                compareStage_counterOnePixelStream_s2mPipe_valid;
  reg                 compareStage_counterOnePixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_counterOnePixelStream_s2mPipe_payload;
  reg                 compareStage_counterOnePixelStream_rValid;
  reg        [7:0]    compareStage_counterOnePixelStream_rData;
  wire                diffStage_counterOnePixelStream_valid;
  wire                diffStage_counterOnePixelStream_ready;
  wire       [7:0]    diffStage_counterOnePixelStream_payload;
  reg                 compareStage_counterOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_counterOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_42;
  wire                compareStage_mainTwoPixelStream_s2mPipe_valid;
  reg                 compareStage_mainTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_mainTwoPixelStream_s2mPipe_payload;
  reg                 compareStage_mainTwoPixelStream_rValid;
  reg        [7:0]    compareStage_mainTwoPixelStream_rData;
  wire                diffStage_mainTwoPixelStream_valid;
  wire                diffStage_mainTwoPixelStream_ready;
  wire       [7:0]    diffStage_mainTwoPixelStream_payload;
  reg                 compareStage_mainTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_mainTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_43;
  wire                compareStage_counterTwoPixelStream_s2mPipe_valid;
  reg                 compareStage_counterTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_counterTwoPixelStream_s2mPipe_payload;
  reg                 compareStage_counterTwoPixelStream_rValid;
  reg        [7:0]    compareStage_counterTwoPixelStream_rData;
  wire                diffStage_counterTwoPixelStream_valid;
  wire                diffStage_counterTwoPixelStream_ready;
  wire       [7:0]    diffStage_counterTwoPixelStream_payload;
  reg                 compareStage_counterTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_counterTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_44;
  wire                compareStage_mainThreePixelStream_s2mPipe_valid;
  reg                 compareStage_mainThreePixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_mainThreePixelStream_s2mPipe_payload;
  reg                 compareStage_mainThreePixelStream_rValid;
  reg        [7:0]    compareStage_mainThreePixelStream_rData;
  wire                diffStage_mainThreePixelStream_valid;
  wire                diffStage_mainThreePixelStream_ready;
  wire       [7:0]    diffStage_mainThreePixelStream_payload;
  reg                 compareStage_mainThreePixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_mainThreePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_45;
  wire                compareStage_counterThreePixelStream_s2mPipe_valid;
  reg                 compareStage_counterThreePixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_counterThreePixelStream_s2mPipe_payload;
  reg                 compareStage_counterThreePixelStream_rValid;
  reg        [7:0]    compareStage_counterThreePixelStream_rData;
  wire                diffStage_counterThreePixelStream_valid;
  wire                diffStage_counterThreePixelStream_ready;
  wire       [7:0]    diffStage_counterThreePixelStream_payload;
  reg                 compareStage_counterThreePixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_counterThreePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_46;
  wire                compareStage_mainOneValidStream_s2mPipe_valid;
  reg                 compareStage_mainOneValidStream_s2mPipe_ready;
  wire                compareStage_mainOneValidStream_s2mPipe_payload;
  reg                 compareStage_mainOneValidStream_rValid;
  reg                 compareStage_mainOneValidStream_rData;
  wire                diffStage_mainOneValidStream_valid;
  wire                diffStage_mainOneValidStream_ready;
  wire                diffStage_mainOneValidStream_payload;
  reg                 compareStage_mainOneValidStream_s2mPipe_rValid;
  reg                 compareStage_mainOneValidStream_s2mPipe_rData;
  wire                when_Stream_l368_47;
  wire                compareStage_counterOneValidStream_s2mPipe_valid;
  reg                 compareStage_counterOneValidStream_s2mPipe_ready;
  wire                compareStage_counterOneValidStream_s2mPipe_payload;
  reg                 compareStage_counterOneValidStream_rValid;
  reg                 compareStage_counterOneValidStream_rData;
  wire                diffStage_counterOneValidStream_valid;
  wire                diffStage_counterOneValidStream_ready;
  wire                diffStage_counterOneValidStream_payload;
  reg                 compareStage_counterOneValidStream_s2mPipe_rValid;
  reg                 compareStage_counterOneValidStream_s2mPipe_rData;
  wire                when_Stream_l368_48;
  wire                compareStage_mainTwoValidStream_s2mPipe_valid;
  reg                 compareStage_mainTwoValidStream_s2mPipe_ready;
  wire                compareStage_mainTwoValidStream_s2mPipe_payload;
  reg                 compareStage_mainTwoValidStream_rValid;
  reg                 compareStage_mainTwoValidStream_rData;
  wire                diffStage_mainTwoValidStream_valid;
  wire                diffStage_mainTwoValidStream_ready;
  wire                diffStage_mainTwoValidStream_payload;
  reg                 compareStage_mainTwoValidStream_s2mPipe_rValid;
  reg                 compareStage_mainTwoValidStream_s2mPipe_rData;
  wire                when_Stream_l368_49;
  wire                compareStage_counterTwoValidStream_s2mPipe_valid;
  reg                 compareStage_counterTwoValidStream_s2mPipe_ready;
  wire                compareStage_counterTwoValidStream_s2mPipe_payload;
  reg                 compareStage_counterTwoValidStream_rValid;
  reg                 compareStage_counterTwoValidStream_rData;
  wire                diffStage_counterTwoValidStream_valid;
  wire                diffStage_counterTwoValidStream_ready;
  wire                diffStage_counterTwoValidStream_payload;
  reg                 compareStage_counterTwoValidStream_s2mPipe_rValid;
  reg                 compareStage_counterTwoValidStream_s2mPipe_rData;
  wire                when_Stream_l368_50;
  wire                compareStage_mainThreeValidStream_s2mPipe_valid;
  reg                 compareStage_mainThreeValidStream_s2mPipe_ready;
  wire                compareStage_mainThreeValidStream_s2mPipe_payload;
  reg                 compareStage_mainThreeValidStream_rValid;
  reg                 compareStage_mainThreeValidStream_rData;
  wire                diffStage_mainThreeValidStream_valid;
  wire                diffStage_mainThreeValidStream_ready;
  wire                diffStage_mainThreeValidStream_payload;
  reg                 compareStage_mainThreeValidStream_s2mPipe_rValid;
  reg                 compareStage_mainThreeValidStream_s2mPipe_rData;
  wire                when_Stream_l368_51;
  wire                compareStage_counterThreeValidStream_s2mPipe_valid;
  reg                 compareStage_counterThreeValidStream_s2mPipe_ready;
  wire                compareStage_counterThreeValidStream_s2mPipe_payload;
  reg                 compareStage_counterThreeValidStream_rValid;
  reg                 compareStage_counterThreeValidStream_rData;
  wire                diffStage_counterThreeValidStream_valid;
  wire                diffStage_counterThreeValidStream_ready;
  wire                diffStage_counterThreeValidStream_payload;
  reg                 compareStage_counterThreeValidStream_s2mPipe_rValid;
  reg                 compareStage_counterThreeValidStream_s2mPipe_rData;
  wire                when_Stream_l368_52;
  reg        [7:0]    CICC1851_compareStage_controlPipe_translated_payload_mainDiff;
  reg        [7:0]    CICC1851_compareStage_controlPipe_translated_payload_counterDiff;
  reg        [7:0]    CICC1851_compareStage_controlPipe_translated_payload_horizontalDiff;
  reg        [7:0]    CICC1851_compareStage_controlPipe_translated_payload_verticalDiff;
  reg                 CICC1851_compareStage_controlPipe_translated_payload_inValidMinDiff;
  wire                when_SuperResolutionPart3_l647;
  wire                when_SuperResolutionPart3_l649;
  wire                when_SuperResolutionPart3_l652;
  wire                when_SuperResolutionPart3_l661;
  wire                when_SuperResolutionPart3_l664;
  wire                when_SuperResolutionPart3_l697;
  wire                when_SuperResolutionPart3_l725;
  wire                when_SuperResolutionPart3_l694;
  wire                when_SuperResolutionPart3_l753;
  wire                compareStage_controlPipe_translated_valid;
  wire                compareStage_controlPipe_translated_ready;
  wire                compareStage_controlPipe_translated_payload_frameStart;
  wire                compareStage_controlPipe_translated_payload_rowEnd;
  wire                compareStage_controlPipe_translated_payload_pipeValid;
  wire                compareStage_controlPipe_translated_payload_firstRow;
  wire                compareStage_controlPipe_translated_payload_lastRow;
  wire                compareStage_controlPipe_translated_payload_finalResult;
  wire                compareStage_controlPipe_translated_payload_mainCompare;
  wire                compareStage_controlPipe_translated_payload_counterCompare;
  wire                compareStage_controlPipe_translated_payload_horizontalCompare;
  wire                compareStage_controlPipe_translated_payload_verticalCompare;
  wire       [7:0]    compareStage_controlPipe_translated_payload_mainDiff;
  wire       [7:0]    compareStage_controlPipe_translated_payload_counterDiff;
  wire       [7:0]    compareStage_controlPipe_translated_payload_horizontalDiff;
  wire       [7:0]    compareStage_controlPipe_translated_payload_verticalDiff;
  wire                compareStage_controlPipe_translated_payload_isHorizontalMin;
  wire       [7:0]    compareStage_controlPipe_translated_payload_minDiff;
  wire       [1:0]    compareStage_controlPipe_translated_payload_currentPosition;
  wire       [1:0]    compareStage_controlPipe_translated_payload_nextPosition;
  wire                compareStage_controlPipe_translated_payload_horizontalDirectionValid;
  wire                compareStage_controlPipe_translated_payload_verticalDirectionValid;
  wire                compareStage_controlPipe_translated_payload_mainDirectionValid;
  wire                compareStage_controlPipe_translated_payload_counterDirectionValid;
  wire                compareStage_controlPipe_translated_payload_inValidMinDiff;
  wire                compareStage_controlPipe_translated_s2mPipe_valid;
  reg                 compareStage_controlPipe_translated_s2mPipe_ready;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_frameStart;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_rowEnd;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_pipeValid;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_firstRow;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_lastRow;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_finalResult;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_mainCompare;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_counterCompare;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_horizontalCompare;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_verticalCompare;
  wire       [7:0]    compareStage_controlPipe_translated_s2mPipe_payload_mainDiff;
  wire       [7:0]    compareStage_controlPipe_translated_s2mPipe_payload_counterDiff;
  wire       [7:0]    compareStage_controlPipe_translated_s2mPipe_payload_horizontalDiff;
  wire       [7:0]    compareStage_controlPipe_translated_s2mPipe_payload_verticalDiff;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_isHorizontalMin;
  wire       [7:0]    compareStage_controlPipe_translated_s2mPipe_payload_minDiff;
  wire       [1:0]    compareStage_controlPipe_translated_s2mPipe_payload_currentPosition;
  wire       [1:0]    compareStage_controlPipe_translated_s2mPipe_payload_nextPosition;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_horizontalDirectionValid;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_verticalDirectionValid;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_mainDirectionValid;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_counterDirectionValid;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_inValidMinDiff;
  reg                 compareStage_controlPipe_translated_rValid;
  reg                 compareStage_controlPipe_translated_rData_frameStart;
  reg                 compareStage_controlPipe_translated_rData_rowEnd;
  reg                 compareStage_controlPipe_translated_rData_pipeValid;
  reg                 compareStage_controlPipe_translated_rData_firstRow;
  reg                 compareStage_controlPipe_translated_rData_lastRow;
  reg                 compareStage_controlPipe_translated_rData_finalResult;
  reg                 compareStage_controlPipe_translated_rData_mainCompare;
  reg                 compareStage_controlPipe_translated_rData_counterCompare;
  reg                 compareStage_controlPipe_translated_rData_horizontalCompare;
  reg                 compareStage_controlPipe_translated_rData_verticalCompare;
  reg        [7:0]    compareStage_controlPipe_translated_rData_mainDiff;
  reg        [7:0]    compareStage_controlPipe_translated_rData_counterDiff;
  reg        [7:0]    compareStage_controlPipe_translated_rData_horizontalDiff;
  reg        [7:0]    compareStage_controlPipe_translated_rData_verticalDiff;
  reg                 compareStage_controlPipe_translated_rData_isHorizontalMin;
  reg        [7:0]    compareStage_controlPipe_translated_rData_minDiff;
  reg        [1:0]    compareStage_controlPipe_translated_rData_currentPosition;
  reg        [1:0]    compareStage_controlPipe_translated_rData_nextPosition;
  reg                 compareStage_controlPipe_translated_rData_horizontalDirectionValid;
  reg                 compareStage_controlPipe_translated_rData_verticalDirectionValid;
  reg                 compareStage_controlPipe_translated_rData_mainDirectionValid;
  reg                 compareStage_controlPipe_translated_rData_counterDirectionValid;
  reg                 compareStage_controlPipe_translated_rData_inValidMinDiff;
  wire                diffStage_controlPipe_valid;
  wire                diffStage_controlPipe_ready;
  wire                diffStage_controlPipe_payload_frameStart;
  wire                diffStage_controlPipe_payload_rowEnd;
  wire                diffStage_controlPipe_payload_pipeValid;
  wire                diffStage_controlPipe_payload_firstRow;
  wire                diffStage_controlPipe_payload_lastRow;
  wire                diffStage_controlPipe_payload_finalResult;
  wire                diffStage_controlPipe_payload_mainCompare;
  wire                diffStage_controlPipe_payload_counterCompare;
  wire                diffStage_controlPipe_payload_horizontalCompare;
  wire                diffStage_controlPipe_payload_verticalCompare;
  wire       [7:0]    diffStage_controlPipe_payload_mainDiff;
  wire       [7:0]    diffStage_controlPipe_payload_counterDiff;
  wire       [7:0]    diffStage_controlPipe_payload_horizontalDiff;
  wire       [7:0]    diffStage_controlPipe_payload_verticalDiff;
  wire                diffStage_controlPipe_payload_isHorizontalMin;
  wire       [7:0]    diffStage_controlPipe_payload_minDiff;
  wire       [1:0]    diffStage_controlPipe_payload_currentPosition;
  wire       [1:0]    diffStage_controlPipe_payload_nextPosition;
  wire                diffStage_controlPipe_payload_horizontalDirectionValid;
  wire                diffStage_controlPipe_payload_verticalDirectionValid;
  wire                diffStage_controlPipe_payload_mainDirectionValid;
  wire                diffStage_controlPipe_payload_counterDirectionValid;
  wire                diffStage_controlPipe_payload_inValidMinDiff;
  reg                 compareStage_controlPipe_translated_s2mPipe_rValid;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_frameStart;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_rowEnd;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_pipeValid;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_firstRow;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_lastRow;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_finalResult;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_mainCompare;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_counterCompare;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_horizontalCompare;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_verticalCompare;
  reg        [7:0]    compareStage_controlPipe_translated_s2mPipe_rData_mainDiff;
  reg        [7:0]    compareStage_controlPipe_translated_s2mPipe_rData_counterDiff;
  reg        [7:0]    compareStage_controlPipe_translated_s2mPipe_rData_horizontalDiff;
  reg        [7:0]    compareStage_controlPipe_translated_s2mPipe_rData_verticalDiff;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_isHorizontalMin;
  reg        [7:0]    compareStage_controlPipe_translated_s2mPipe_rData_minDiff;
  reg        [1:0]    compareStage_controlPipe_translated_s2mPipe_rData_currentPosition;
  reg        [1:0]    compareStage_controlPipe_translated_s2mPipe_rData_nextPosition;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_horizontalDirectionValid;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_verticalDirectionValid;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_mainDirectionValid;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_counterDirectionValid;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_inValidMinDiff;
  wire                when_Stream_l368_53;
  wire                diffStage_mainOnePixelStream_s2mPipe_valid;
  reg                 diffStage_mainOnePixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_mainOnePixelStream_s2mPipe_payload;
  reg                 diffStage_mainOnePixelStream_rValid;
  reg        [7:0]    diffStage_mainOnePixelStream_rData;
  wire                resultStage_mainOnePixelStream_valid;
  wire                resultStage_mainOnePixelStream_ready;
  wire       [7:0]    resultStage_mainOnePixelStream_payload;
  reg                 diffStage_mainOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_mainOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_54;
  wire                diffStage_counterOnePixelStream_s2mPipe_valid;
  reg                 diffStage_counterOnePixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_counterOnePixelStream_s2mPipe_payload;
  reg                 diffStage_counterOnePixelStream_rValid;
  reg        [7:0]    diffStage_counterOnePixelStream_rData;
  wire                resultStage_counterOnePixelStream_valid;
  wire                resultStage_counterOnePixelStream_ready;
  wire       [7:0]    resultStage_counterOnePixelStream_payload;
  reg                 diffStage_counterOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_counterOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_55;
  wire                diffStage_mainTwoPixelStream_s2mPipe_valid;
  reg                 diffStage_mainTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_mainTwoPixelStream_s2mPipe_payload;
  reg                 diffStage_mainTwoPixelStream_rValid;
  reg        [7:0]    diffStage_mainTwoPixelStream_rData;
  wire                resultStage_mainTwoPixelStream_valid;
  wire                resultStage_mainTwoPixelStream_ready;
  wire       [7:0]    resultStage_mainTwoPixelStream_payload;
  reg                 diffStage_mainTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_mainTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_56;
  wire                diffStage_counterTwoPixelStream_s2mPipe_valid;
  reg                 diffStage_counterTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_counterTwoPixelStream_s2mPipe_payload;
  reg                 diffStage_counterTwoPixelStream_rValid;
  reg        [7:0]    diffStage_counterTwoPixelStream_rData;
  wire                resultStage_counterTwoPixelStream_valid;
  wire                resultStage_counterTwoPixelStream_ready;
  wire       [7:0]    resultStage_counterTwoPixelStream_payload;
  reg                 diffStage_counterTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_counterTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_57;
  wire                diffStage_mainThreePixelStream_s2mPipe_valid;
  reg                 diffStage_mainThreePixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_mainThreePixelStream_s2mPipe_payload;
  reg                 diffStage_mainThreePixelStream_rValid;
  reg        [7:0]    diffStage_mainThreePixelStream_rData;
  wire                resultStage_mainThreePixelStream_valid;
  wire                resultStage_mainThreePixelStream_ready;
  wire       [7:0]    resultStage_mainThreePixelStream_payload;
  reg                 diffStage_mainThreePixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_mainThreePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_58;
  wire                diffStage_counterThreePixelStream_s2mPipe_valid;
  reg                 diffStage_counterThreePixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_counterThreePixelStream_s2mPipe_payload;
  reg                 diffStage_counterThreePixelStream_rValid;
  reg        [7:0]    diffStage_counterThreePixelStream_rData;
  wire                resultStage_counterThreePixelStream_valid;
  wire                resultStage_counterThreePixelStream_ready;
  wire       [7:0]    resultStage_counterThreePixelStream_payload;
  reg                 diffStage_counterThreePixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_counterThreePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_59;
  wire                diffStage_mainOneValidStream_s2mPipe_valid;
  reg                 diffStage_mainOneValidStream_s2mPipe_ready;
  wire                diffStage_mainOneValidStream_s2mPipe_payload;
  reg                 diffStage_mainOneValidStream_rValid;
  reg                 diffStage_mainOneValidStream_rData;
  wire                resultStage_mainOneValidStream_valid;
  wire                resultStage_mainOneValidStream_ready;
  wire                resultStage_mainOneValidStream_payload;
  reg                 diffStage_mainOneValidStream_s2mPipe_rValid;
  reg                 diffStage_mainOneValidStream_s2mPipe_rData;
  wire                when_Stream_l368_60;
  wire                diffStage_counterOneValidStream_s2mPipe_valid;
  reg                 diffStage_counterOneValidStream_s2mPipe_ready;
  wire                diffStage_counterOneValidStream_s2mPipe_payload;
  reg                 diffStage_counterOneValidStream_rValid;
  reg                 diffStage_counterOneValidStream_rData;
  wire                resultStage_counterOneValidStream_valid;
  wire                resultStage_counterOneValidStream_ready;
  wire                resultStage_counterOneValidStream_payload;
  reg                 diffStage_counterOneValidStream_s2mPipe_rValid;
  reg                 diffStage_counterOneValidStream_s2mPipe_rData;
  wire                when_Stream_l368_61;
  wire                diffStage_mainTwoValidStream_s2mPipe_valid;
  reg                 diffStage_mainTwoValidStream_s2mPipe_ready;
  wire                diffStage_mainTwoValidStream_s2mPipe_payload;
  reg                 diffStage_mainTwoValidStream_rValid;
  reg                 diffStage_mainTwoValidStream_rData;
  wire                resultStage_mainTwoValidStream_valid;
  wire                resultStage_mainTwoValidStream_ready;
  wire                resultStage_mainTwoValidStream_payload;
  reg                 diffStage_mainTwoValidStream_s2mPipe_rValid;
  reg                 diffStage_mainTwoValidStream_s2mPipe_rData;
  wire                when_Stream_l368_62;
  wire                diffStage_counterTwoValidStream_s2mPipe_valid;
  reg                 diffStage_counterTwoValidStream_s2mPipe_ready;
  wire                diffStage_counterTwoValidStream_s2mPipe_payload;
  reg                 diffStage_counterTwoValidStream_rValid;
  reg                 diffStage_counterTwoValidStream_rData;
  wire                resultStage_counterTwoValidStream_valid;
  wire                resultStage_counterTwoValidStream_ready;
  wire                resultStage_counterTwoValidStream_payload;
  reg                 diffStage_counterTwoValidStream_s2mPipe_rValid;
  reg                 diffStage_counterTwoValidStream_s2mPipe_rData;
  wire                when_Stream_l368_63;
  wire                diffStage_mainThreeValidStream_s2mPipe_valid;
  reg                 diffStage_mainThreeValidStream_s2mPipe_ready;
  wire                diffStage_mainThreeValidStream_s2mPipe_payload;
  reg                 diffStage_mainThreeValidStream_rValid;
  reg                 diffStage_mainThreeValidStream_rData;
  wire                resultStage_mainThreeValidStream_valid;
  wire                resultStage_mainThreeValidStream_ready;
  wire                resultStage_mainThreeValidStream_payload;
  reg                 diffStage_mainThreeValidStream_s2mPipe_rValid;
  reg                 diffStage_mainThreeValidStream_s2mPipe_rData;
  wire                when_Stream_l368_64;
  wire                diffStage_counterThreeValidStream_s2mPipe_valid;
  reg                 diffStage_counterThreeValidStream_s2mPipe_ready;
  wire                diffStage_counterThreeValidStream_s2mPipe_payload;
  reg                 diffStage_counterThreeValidStream_rValid;
  reg                 diffStage_counterThreeValidStream_rData;
  wire                resultStage_counterThreeValidStream_valid;
  wire                resultStage_counterThreeValidStream_ready;
  wire                resultStage_counterThreeValidStream_payload;
  reg                 diffStage_counterThreeValidStream_s2mPipe_rValid;
  reg                 diffStage_counterThreeValidStream_s2mPipe_rData;
  wire                when_Stream_l368_65;
  reg                 CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin;
  reg        [7:0]    CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff;
  wire                when_SuperResolutionPart3_l783;
  wire                when_SuperResolutionPart3_l784;
  wire                when_SuperResolutionPart3_l785;
  wire                when_SuperResolutionPart3_l788;
  wire                when_SuperResolutionPart3_l796;
  wire                when_SuperResolutionPart3_l804;
  wire                when_SuperResolutionPart3_l812;
  wire                when_SuperResolutionPart3_l795;
  wire                when_SuperResolutionPart3_l803;
  wire                when_SuperResolutionPart3_l811;
  wire                when_SuperResolutionPart3_l819;
  wire                when_SuperResolutionPart3_l822;
  wire                when_SuperResolutionPart3_l825;
  wire                resultStage_controlPipeBeforePipe_valid;
  wire                resultStage_controlPipeBeforePipe_ready;
  wire                resultStage_controlPipeBeforePipe_payload_frameStart;
  wire                resultStage_controlPipeBeforePipe_payload_rowEnd;
  wire                resultStage_controlPipeBeforePipe_payload_pipeValid;
  wire                resultStage_controlPipeBeforePipe_payload_firstRow;
  wire                resultStage_controlPipeBeforePipe_payload_lastRow;
  wire                resultStage_controlPipeBeforePipe_payload_finalResult;
  wire                resultStage_controlPipeBeforePipe_payload_mainCompare;
  wire                resultStage_controlPipeBeforePipe_payload_counterCompare;
  wire                resultStage_controlPipeBeforePipe_payload_horizontalCompare;
  wire                resultStage_controlPipeBeforePipe_payload_verticalCompare;
  wire       [7:0]    resultStage_controlPipeBeforePipe_payload_mainDiff;
  wire       [7:0]    resultStage_controlPipeBeforePipe_payload_counterDiff;
  wire       [7:0]    resultStage_controlPipeBeforePipe_payload_horizontalDiff;
  wire       [7:0]    resultStage_controlPipeBeforePipe_payload_verticalDiff;
  wire                resultStage_controlPipeBeforePipe_payload_isHorizontalMin;
  wire       [7:0]    resultStage_controlPipeBeforePipe_payload_minDiff;
  wire       [1:0]    resultStage_controlPipeBeforePipe_payload_currentPosition;
  wire       [1:0]    resultStage_controlPipeBeforePipe_payload_nextPosition;
  wire                resultStage_controlPipeBeforePipe_payload_horizontalDirectionValid;
  wire                resultStage_controlPipeBeforePipe_payload_verticalDirectionValid;
  wire                resultStage_controlPipeBeforePipe_payload_mainDirectionValid;
  wire                resultStage_controlPipeBeforePipe_payload_counterDirectionValid;
  wire                resultStage_controlPipeBeforePipe_payload_inValidMinDiff;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_valid;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_ready;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_frameStart;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_rowEnd;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_pipeValid;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_firstRow;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_lastRow;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_finalResult;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_mainCompare;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_counterCompare;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_horizontalCompare;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_verticalCompare;
  wire       [7:0]    resultStage_controlPipeBeforePipe_s2mPipe_payload_mainDiff;
  wire       [7:0]    resultStage_controlPipeBeforePipe_s2mPipe_payload_counterDiff;
  wire       [7:0]    resultStage_controlPipeBeforePipe_s2mPipe_payload_horizontalDiff;
  wire       [7:0]    resultStage_controlPipeBeforePipe_s2mPipe_payload_verticalDiff;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_isHorizontalMin;
  wire       [7:0]    resultStage_controlPipeBeforePipe_s2mPipe_payload_minDiff;
  wire       [1:0]    resultStage_controlPipeBeforePipe_s2mPipe_payload_currentPosition;
  wire       [1:0]    resultStage_controlPipeBeforePipe_s2mPipe_payload_nextPosition;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_horizontalDirectionValid;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_verticalDirectionValid;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_mainDirectionValid;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_counterDirectionValid;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_inValidMinDiff;
  reg                 resultStage_controlPipeBeforePipe_rValid;
  reg                 resultStage_controlPipeBeforePipe_rData_frameStart;
  reg                 resultStage_controlPipeBeforePipe_rData_rowEnd;
  reg                 resultStage_controlPipeBeforePipe_rData_pipeValid;
  reg                 resultStage_controlPipeBeforePipe_rData_firstRow;
  reg                 resultStage_controlPipeBeforePipe_rData_lastRow;
  reg                 resultStage_controlPipeBeforePipe_rData_finalResult;
  reg                 resultStage_controlPipeBeforePipe_rData_mainCompare;
  reg                 resultStage_controlPipeBeforePipe_rData_counterCompare;
  reg                 resultStage_controlPipeBeforePipe_rData_horizontalCompare;
  reg                 resultStage_controlPipeBeforePipe_rData_verticalCompare;
  reg        [7:0]    resultStage_controlPipeBeforePipe_rData_mainDiff;
  reg        [7:0]    resultStage_controlPipeBeforePipe_rData_counterDiff;
  reg        [7:0]    resultStage_controlPipeBeforePipe_rData_horizontalDiff;
  reg        [7:0]    resultStage_controlPipeBeforePipe_rData_verticalDiff;
  reg                 resultStage_controlPipeBeforePipe_rData_isHorizontalMin;
  reg        [7:0]    resultStage_controlPipeBeforePipe_rData_minDiff;
  reg        [1:0]    resultStage_controlPipeBeforePipe_rData_currentPosition;
  reg        [1:0]    resultStage_controlPipeBeforePipe_rData_nextPosition;
  reg                 resultStage_controlPipeBeforePipe_rData_horizontalDirectionValid;
  reg                 resultStage_controlPipeBeforePipe_rData_verticalDirectionValid;
  reg                 resultStage_controlPipeBeforePipe_rData_mainDirectionValid;
  reg                 resultStage_controlPipeBeforePipe_rData_counterDirectionValid;
  reg                 resultStage_controlPipeBeforePipe_rData_inValidMinDiff;
  wire                resultStage_controlPipe_valid;
  wire                resultStage_controlPipe_ready;
  wire                resultStage_controlPipe_payload_frameStart;
  wire                resultStage_controlPipe_payload_rowEnd;
  wire                resultStage_controlPipe_payload_pipeValid;
  wire                resultStage_controlPipe_payload_firstRow;
  wire                resultStage_controlPipe_payload_lastRow;
  wire                resultStage_controlPipe_payload_finalResult;
  wire                resultStage_controlPipe_payload_mainCompare;
  wire                resultStage_controlPipe_payload_counterCompare;
  wire                resultStage_controlPipe_payload_horizontalCompare;
  wire                resultStage_controlPipe_payload_verticalCompare;
  wire       [7:0]    resultStage_controlPipe_payload_mainDiff;
  wire       [7:0]    resultStage_controlPipe_payload_counterDiff;
  wire       [7:0]    resultStage_controlPipe_payload_horizontalDiff;
  wire       [7:0]    resultStage_controlPipe_payload_verticalDiff;
  wire                resultStage_controlPipe_payload_isHorizontalMin;
  wire       [7:0]    resultStage_controlPipe_payload_minDiff;
  wire       [1:0]    resultStage_controlPipe_payload_currentPosition;
  wire       [1:0]    resultStage_controlPipe_payload_nextPosition;
  wire                resultStage_controlPipe_payload_horizontalDirectionValid;
  wire                resultStage_controlPipe_payload_verticalDirectionValid;
  wire                resultStage_controlPipe_payload_mainDirectionValid;
  wire                resultStage_controlPipe_payload_counterDirectionValid;
  wire                resultStage_controlPipe_payload_inValidMinDiff;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rValid;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_frameStart;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_rowEnd;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_pipeValid;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_firstRow;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_lastRow;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_finalResult;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_mainCompare;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_counterCompare;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_horizontalCompare;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_verticalCompare;
  reg        [7:0]    resultStage_controlPipeBeforePipe_s2mPipe_rData_mainDiff;
  reg        [7:0]    resultStage_controlPipeBeforePipe_s2mPipe_rData_counterDiff;
  reg        [7:0]    resultStage_controlPipeBeforePipe_s2mPipe_rData_horizontalDiff;
  reg        [7:0]    resultStage_controlPipeBeforePipe_s2mPipe_rData_verticalDiff;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_isHorizontalMin;
  reg        [7:0]    resultStage_controlPipeBeforePipe_s2mPipe_rData_minDiff;
  reg        [1:0]    resultStage_controlPipeBeforePipe_s2mPipe_rData_currentPosition;
  reg        [1:0]    resultStage_controlPipeBeforePipe_s2mPipe_rData_nextPosition;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_horizontalDirectionValid;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_verticalDirectionValid;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_mainDirectionValid;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_counterDirectionValid;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_inValidMinDiff;
  wire                when_Stream_l368_66;
  wire                resultStage_pixelStream_valid;
  wire                resultStage_pixelStream_ready;
  reg        [7:0]    resultStage_pixelStream_payload;
  wire                when_SuperResolutionPart3_l840;
  wire                when_SuperResolutionPart3_l846;
  wire                when_SuperResolutionPart3_l847;
  wire                when_SuperResolutionPart3_l850;
  wire                when_SuperResolutionPart3_l854;
  wire                when_SuperResolutionPart3_l855;
  wire                when_SuperResolutionPart3_l860;
  wire                when_SuperResolutionPart3_l861;
  wire                when_SuperResolutionPart3_l851;
  wire                when_SuperResolutionPart3_l841;
  wire                when_SuperResolutionPart3_l842;
  wire                when_SuperResolutionPart3_l869;
  wire                when_SuperResolutionPart3_l870;
  wire                when_SuperResolutionPart3_l871;
  wire                when_SuperResolutionPart3_l872;
  wire                when_SuperResolutionPart3_l875;
  wire                when_SuperResolutionPart3_l876;
  wire                when_SuperResolutionPart3_l885;
  wire                when_SuperResolutionPart3_l893;
  wire                when_SuperResolutionPart3_l884;
  wire                when_SuperResolutionPart3_l902;
  wire                when_SuperResolutionPart3_l903;
  wire                when_SuperResolutionPart3_l912;
  wire                when_SuperResolutionPart3_l920;
  wire                when_SuperResolutionPart3_l911;
  wire                when_SuperResolutionPart3_l874;
  wire                when_SuperResolutionPart3_l930;
  wire                when_SuperResolutionPart3_l931;
  wire                when_SuperResolutionPart3_l932;
  wire                when_SuperResolutionPart3_l941;
  wire                when_SuperResolutionPart3_l949;
  wire                when_SuperResolutionPart3_l940;
  wire                when_SuperResolutionPart3_l958;
  wire                when_SuperResolutionPart3_l959;
  wire                when_SuperResolutionPart3_l968;
  wire                when_SuperResolutionPart3_l976;
  wire                when_SuperResolutionPart3_l967;
  wire                when_SuperResolutionPart3_l986;
  wire                when_SuperResolutionPart3_l987;
  wire                when_SuperResolutionPart3_l988;
  wire                when_SuperResolutionPart3_l991;
  wire                when_SuperResolutionPart3_l992;
  wire                when_SuperResolutionPart3_l1001;
  wire                when_SuperResolutionPart3_l1009;
  wire                when_SuperResolutionPart3_l1000;
  wire                when_SuperResolutionPart3_l1019;
  wire                when_SuperResolutionPart3_l1020;
  wire                when_SuperResolutionPart3_l1021;
  wire                when_SuperResolutionPart3_l1024;
  wire                when_SuperResolutionPart3_l1025;
  wire                when_SuperResolutionPart3_l1034;
  wire                when_SuperResolutionPart3_l1042;
  wire                when_SuperResolutionPart3_l1033;
  wire                when_SuperResolutionPart3_l1052;
  wire                when_SuperResolutionPart3_l1053;
  wire                when_SuperResolutionPart3_l1062;
  wire                when_SuperResolutionPart3_l1070;
  wire                when_SuperResolutionPart3_l1061;
  wire                when_SuperResolutionPart3_l1079;
  wire                when_SuperResolutionPart3_l1080;
  wire                when_SuperResolutionPart3_l1083;
  wire                when_SuperResolutionPart3_l1084;
  wire                when_SuperResolutionPart3_l1093;
  wire                when_SuperResolutionPart3_l1101;
  wire                when_SuperResolutionPart3_l1092;
  wire                when_SuperResolutionPart3_l929;
  wire                when_SuperResolutionPart3_l985;
  wire                when_SuperResolutionPart3_l1018;
  wire                when_SuperResolutionPart3_l1051;
  wire                when_SuperResolutionPart3_l1078;
  wire                when_SuperResolutionPart3_l1082;
  wire                resultStage_pixelStream_s2mPipe_valid;
  reg                 resultStage_pixelStream_s2mPipe_ready;
  wire       [7:0]    resultStage_pixelStream_s2mPipe_payload;
  reg                 resultStage_pixelStream_rValid;
  reg        [7:0]    resultStage_pixelStream_rData;
  wire                resultStage_resultStream_valid;
  wire                resultStage_resultStream_ready;
  wire       [7:0]    resultStage_resultStream_payload;
  reg                 resultStage_pixelStream_s2mPipe_rValid;
  reg        [7:0]    resultStage_pixelStream_s2mPipe_rData;
  wire                when_Stream_l368_67;
  wire                when_SuperResolutionPart3_l1115;
  wire                diffStage_controlPipe_fire;
  wire                CICC1851_resultStage_mainOnePixelStream_ready;
  reg                 CICC1851_resultStage_mainOnePixelStream_ready_1;
  wire                CICC1851_resultStage_mainOnePixelStream_ready_2;
  wire                when_Stream_l438;
  reg                 resultsJoin_valid;
  wire                resultsJoin_ready;
  wire                pixelsStream_valid;
  wire                pixelsStream_ready;
  wire       [7:0]    pixelsStream_payload_pixel;
  wire                pixelsStream_payload_frameStart;
  wire                pixelsStream_payload_rowEnd;
  wire                pixelsStream_s2mPipe_valid;
  reg                 pixelsStream_s2mPipe_ready;
  wire       [7:0]    pixelsStream_s2mPipe_payload_pixel;
  wire                pixelsStream_s2mPipe_payload_frameStart;
  wire                pixelsStream_s2mPipe_payload_rowEnd;
  reg                 pixelsStream_rValid;
  reg        [7:0]    pixelsStream_rData_pixel;
  reg                 pixelsStream_rData_frameStart;
  reg                 pixelsStream_rData_rowEnd;
  wire                pixelsStream_s2mPipe_m2sPipe_valid;
  wire                pixelsStream_s2mPipe_m2sPipe_ready;
  wire       [7:0]    pixelsStream_s2mPipe_m2sPipe_payload_pixel;
  wire                pixelsStream_s2mPipe_m2sPipe_payload_frameStart;
  wire                pixelsStream_s2mPipe_m2sPipe_payload_rowEnd;
  reg                 pixelsStream_s2mPipe_rValid;
  reg        [7:0]    pixelsStream_s2mPipe_rData_pixel;
  reg                 pixelsStream_s2mPipe_rData_frameStart;
  reg                 pixelsStream_s2mPipe_rData_rowEnd;
  wire                when_Stream_l368_68;
  wire                controlStateMachine_wantExit;
  reg                 controlStateMachine_wantStart;
  wire                controlStateMachine_wantKill;
  reg        [1:0]    controlStateMachine_stateReg;
  reg        [1:0]    controlStateMachine_stateNext;
  wire                passPixels_fire_13;
  wire                when_SuperResolutionPart3_l1158;
  wire                controlStream_fire;
  wire                when_SuperResolutionPart3_l1168;
  wire                when_SuperResolutionPart3_l1188;
  wire                controlStream_fire_1;
  wire                when_SuperResolutionPart3_l1199;
  wire                passPixels_fire_14;
  wire                when_SuperResolutionPart3_l1202;
  wire                passPixels_fire_15;
  wire                when_SuperResolutionPart3_l1205;
  wire                when_SuperResolutionPart3_l1217;
  wire                controlStream_fire_2;
  wire                when_SuperResolutionPart3_l1220;
  wire                controlStream_fire_3;
  wire                when_SuperResolutionPart3_l1223;
  wire                controlStream_fire_4;
  wire                when_SuperResolutionPart3_l1224;
  wire                controlStream_fire_5;
  wire                when_SuperResolutionPart3_l1226;
  wire                controlStream_fire_6;
  wire                controlStream_fire_7;
  wire                when_SuperResolutionPart3_l1247;
  wire                when_SuperResolutionPart3_l1248;
  wire                when_SuperResolutionPart3_l1250;
  wire                when_SuperResolutionPart3_l1252;
  `ifndef SYNTHESIS
  reg [39:0] controlStateMachine_stateReg_string;
  reg [39:0] controlStateMachine_stateNext_string;
  `endif

  reg [7:0] lineBufferOne [0:3839];
  reg [7:0] lineBufferTwo [0:3839];
  reg [7:0] lineBufferThree [0:3839];
  reg [0:0] validBufferOne [0:3839];
  reg [0:0] validBufferTwo [0:3839];
  reg [0:0] validBufferThree [0:3839];

  assign CICC1851_bufferRowCount_valueNext_1 = bufferRowCount_willIncrement;
  assign CICC1851_bufferRowCount_valueNext = {11'd0, CICC1851_bufferRowCount_valueNext_1};
  assign CICC1851_bufferWAddr_valueNext_1 = bufferWAddr_willIncrement;
  assign CICC1851_bufferWAddr_valueNext = {11'd0, CICC1851_bufferWAddr_valueNext_1};
  assign CICC1851_outPixelAddr_valueNext_1 = outPixelAddr_willIncrement;
  assign CICC1851_outPixelAddr_valueNext = {11'd0, CICC1851_outPixelAddr_valueNext_1};
  assign CICC1851_outRowCount_valueNext_1 = outRowCount_willIncrement;
  assign CICC1851_outRowCount_valueNext = {11'd0, CICC1851_outRowCount_valueNext_1};
  assign CICC1851_alreadySendRow_valueNext_1 = alreadySendRow_willIncrement;
  assign CICC1851_alreadySendRow_valueNext = {11'd0, CICC1851_alreadySendRow_valueNext_1};
  assign CICC1851_alreadySendCountInRow_valueNext_1 = alreadySendCountInRow_willIncrement;
  assign CICC1851_alreadySendCountInRow_valueNext = {11'd0, CICC1851_alreadySendCountInRow_valueNext_1};
  assign CICC1851_nextRowBuffer = 1'b1;
  assign CICC1851_when_SuperResolutionPart3_l226 = {1'd0, bufferWAddr_value};
  assign CICC1851_when_SuperResolutionPart3_l226_1 = (CICC1851_when_SuperResolutionPart3_l226_2 - 13'h0002);
  assign CICC1851_when_SuperResolutionPart3_l226_2 = (3'b100 * bmpWidth);
  assign CICC1851_when_SuperResolutionPart3_l227 = {1'd0, bufferRowCount_value};
  assign CICC1851_when_SuperResolutionPart3_l227_1 = (CICC1851_when_SuperResolutionPart3_l227_2 - 13'h0002);
  assign CICC1851_when_SuperResolutionPart3_l227_2 = (3'b100 * bmpHeight);
  assign CICC1851_when_SuperResolutionPart3_l270 = {1'd0, alreadySendCountInRow_value};
  assign CICC1851_when_SuperResolutionPart3_l270_1 = (CICC1851_when_SuperResolutionPart3_l270_2 - 13'h0002);
  assign CICC1851_when_SuperResolutionPart3_l270_2 = (3'b100 * bmpWidth);
  assign CICC1851_when_SuperResolutionPart3_l271 = {1'd0, alreadySendRow_value};
  assign CICC1851_when_SuperResolutionPart3_l271_1 = (CICC1851_when_SuperResolutionPart3_l271_2 - 13'h0002);
  assign CICC1851_when_SuperResolutionPart3_l271_2 = (3'b100 * bmpHeight);
  assign CICC1851_resultStage_pixelStream_payload = (CICC1851_resultStage_pixelStream_payload_1 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_1 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_mainThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_2 = (CICC1851_resultStage_pixelStream_payload_3 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_3 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_mainThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_4 = (CICC1851_resultStage_pixelStream_payload_5 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_5 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_mainTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_6 = (CICC1851_resultStage_pixelStream_payload_7 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_7 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_mainThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_8 = (CICC1851_resultStage_pixelStream_payload_9 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_9 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_mainThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_10 = (CICC1851_resultStage_pixelStream_payload_11 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_11 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_mainTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_12 = (CICC1851_resultStage_pixelStream_payload_13 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_13 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_mainThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_14 = (CICC1851_resultStage_pixelStream_payload_15 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_15 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_mainThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_16 = (CICC1851_resultStage_pixelStream_payload_17 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_17 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_mainTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_18 = (CICC1851_resultStage_pixelStream_payload_19 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_19 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_20 = (CICC1851_resultStage_pixelStream_payload_21 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_21 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_22 = (CICC1851_resultStage_pixelStream_payload_23 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_23 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_24 = (CICC1851_resultStage_pixelStream_payload_25 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_25 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_26 = (CICC1851_resultStage_pixelStream_payload_27 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_27 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_28 = (CICC1851_resultStage_pixelStream_payload_29 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_29 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_30 = (CICC1851_resultStage_pixelStream_payload_31 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_31 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_32 = (CICC1851_resultStage_pixelStream_payload_33 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_33 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_34 = (CICC1851_resultStage_pixelStream_payload_35 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_35 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_36 = (CICC1851_resultStage_pixelStream_payload_37 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_37 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_38 = (CICC1851_resultStage_pixelStream_payload_39 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_39 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_40 = (CICC1851_resultStage_pixelStream_payload_41 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_41 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_42 = (CICC1851_resultStage_pixelStream_payload_43 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_43 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_44 = (CICC1851_resultStage_pixelStream_payload_45 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_45 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_46 = (CICC1851_resultStage_pixelStream_payload_47 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_47 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_48 = (CICC1851_resultStage_pixelStream_payload_49 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_49 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_50 = (CICC1851_resultStage_pixelStream_payload_51 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_51 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_52 = (CICC1851_resultStage_pixelStream_payload_53 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_53 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_54 = (CICC1851_resultStage_pixelStream_payload_55 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_55 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_56 = (CICC1851_resultStage_pixelStream_payload_57 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_57 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_58 = (CICC1851_resultStage_pixelStream_payload_59 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_59 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_60 = (CICC1851_resultStage_pixelStream_payload_61 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_61 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_62 = (CICC1851_resultStage_pixelStream_payload_63 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_63 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_64 = (CICC1851_resultStage_pixelStream_payload_65 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_65 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_66 = (CICC1851_resultStage_pixelStream_payload_67 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_67 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_68 = (CICC1851_resultStage_pixelStream_payload_69 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_69 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_70 = (CICC1851_resultStage_pixelStream_payload_71 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_71 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_72 = (CICC1851_resultStage_pixelStream_payload_73 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_73 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_74 = (CICC1851_resultStage_pixelStream_payload_75 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_75 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_76 = (CICC1851_resultStage_pixelStream_payload_77 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_77 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_78 = (CICC1851_resultStage_pixelStream_payload_79 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_79 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_80 = (CICC1851_resultStage_pixelStream_payload_81 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_81 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_82 = (CICC1851_resultStage_pixelStream_payload_83 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_83 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_84 = (CICC1851_resultStage_pixelStream_payload_85 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_85 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_86 = (CICC1851_resultStage_pixelStream_payload_87 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_87 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_88 = (CICC1851_resultStage_pixelStream_payload_89 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_89 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_90 = (CICC1851_resultStage_pixelStream_payload_91 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_91 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_92 = (CICC1851_resultStage_pixelStream_payload_93 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_93 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_94 = (CICC1851_resultStage_pixelStream_payload_95 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_95 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_96 = (CICC1851_resultStage_pixelStream_payload_97 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_97 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_98 = (CICC1851_resultStage_pixelStream_payload_99 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_99 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_100 = (CICC1851_resultStage_pixelStream_payload_101 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_101 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_102 = (CICC1851_resultStage_pixelStream_payload_103 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_103 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_104 = (CICC1851_resultStage_pixelStream_payload_105 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_105 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_106 = (CICC1851_resultStage_pixelStream_payload_107 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_107 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_108 = (CICC1851_resultStage_pixelStream_payload_109 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_109 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_110 = (CICC1851_resultStage_pixelStream_payload_111 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_111 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_112 = (CICC1851_resultStage_pixelStream_payload_113 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_113 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_114 = (CICC1851_resultStage_pixelStream_payload_115 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_115 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_116 = (CICC1851_resultStage_pixelStream_payload_117 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_117 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_118 = (CICC1851_resultStage_pixelStream_payload_119 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_119 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_120 = (CICC1851_resultStage_pixelStream_payload_121 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_121 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_122 = (CICC1851_resultStage_pixelStream_payload_123 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_123 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_124 = (CICC1851_resultStage_pixelStream_payload_125 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_125 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_126 = (CICC1851_resultStage_pixelStream_payload_127 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_127 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_128 = (CICC1851_resultStage_pixelStream_payload_129 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_129 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_130 = (CICC1851_resultStage_pixelStream_payload_131 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_131 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_132 = (CICC1851_resultStage_pixelStream_payload_133 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_133 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_134 = (CICC1851_resultStage_pixelStream_payload_135 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_135 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_136 = (CICC1851_resultStage_pixelStream_payload_137 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_137 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_138 = (CICC1851_resultStage_pixelStream_payload_139 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_139 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_140 = (CICC1851_resultStage_pixelStream_payload_141 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_141 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_142 = (CICC1851_resultStage_pixelStream_payload_143 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_143 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_144 = (CICC1851_resultStage_pixelStream_payload_145 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_145 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_146 = (CICC1851_resultStage_pixelStream_payload_147 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_147 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_148 = (CICC1851_resultStage_pixelStream_payload_149 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_149 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_150 = (CICC1851_resultStage_pixelStream_payload_151 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_151 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_152 = (CICC1851_resultStage_pixelStream_payload_153 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_153 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_154 = (CICC1851_resultStage_pixelStream_payload_155 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_155 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_156 = (CICC1851_resultStage_pixelStream_payload_157 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_157 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_158 = (CICC1851_resultStage_pixelStream_payload_159 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_159 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_160 = (CICC1851_resultStage_pixelStream_payload_161 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_161 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_162 = (CICC1851_resultStage_pixelStream_payload_163 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_163 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_164 = (CICC1851_resultStage_pixelStream_payload_165 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_165 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_166 = (CICC1851_resultStage_pixelStream_payload_167 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_167 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_168 = (CICC1851_resultStage_pixelStream_payload_169 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_169 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_170 = (CICC1851_resultStage_pixelStream_payload_171 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_171 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_172 = (CICC1851_resultStage_pixelStream_payload_173 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_173 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_174 = (CICC1851_resultStage_pixelStream_payload_175 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_175 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_176 = (CICC1851_resultStage_pixelStream_payload_177 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_177 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_178 = (CICC1851_resultStage_pixelStream_payload_179 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_179 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_180 = (CICC1851_resultStage_pixelStream_payload_181 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_181 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_182 = (CICC1851_resultStage_pixelStream_payload_183 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_183 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_184 = (CICC1851_resultStage_pixelStream_payload_185 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_185 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_186 = (CICC1851_resultStage_pixelStream_payload_187 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_187 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_188 = (CICC1851_resultStage_pixelStream_payload_189 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_189 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_190 = (CICC1851_resultStage_pixelStream_payload_191 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_191 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_192 = (CICC1851_resultStage_pixelStream_payload_193 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_193 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_194 = (CICC1851_resultStage_pixelStream_payload_195 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_195 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_196 = (CICC1851_resultStage_pixelStream_payload_197 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_197 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_198 = (CICC1851_resultStage_pixelStream_payload_199 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_199 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_200 = (CICC1851_resultStage_pixelStream_payload_201 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_201 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_202 = (CICC1851_resultStage_pixelStream_payload_203 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_203 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_204 = (CICC1851_resultStage_pixelStream_payload_205 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_205 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_206 = (CICC1851_resultStage_pixelStream_payload_207 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_207 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_208 = (CICC1851_resultStage_pixelStream_payload_209 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_209 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_210 = (CICC1851_resultStage_pixelStream_payload_211 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_211 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_212 = (CICC1851_resultStage_pixelStream_payload_213 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_213 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_214 = (CICC1851_resultStage_pixelStream_payload_215 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_215 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_216 = (CICC1851_resultStage_pixelStream_payload_217 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_217 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_218 = (CICC1851_resultStage_pixelStream_payload_219 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_219 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_220 = (CICC1851_resultStage_pixelStream_payload_221 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_221 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_222 = (CICC1851_resultStage_pixelStream_payload_223 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_223 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_224 = (CICC1851_resultStage_pixelStream_payload_225 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_225 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_226 = (CICC1851_resultStage_pixelStream_payload_227 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_227 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_228 = (CICC1851_resultStage_pixelStream_payload_229 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_229 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_230 = (CICC1851_resultStage_pixelStream_payload_231 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_231 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_232 = (CICC1851_resultStage_pixelStream_payload_233 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_233 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_234 = (CICC1851_resultStage_pixelStream_payload_235 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_235 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_236 = (CICC1851_resultStage_pixelStream_payload_237 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_237 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_238 = (CICC1851_resultStage_pixelStream_payload_239 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_239 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_240 = (CICC1851_resultStage_pixelStream_payload_241 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_241 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_242 = (CICC1851_resultStage_pixelStream_payload_243 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_243 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_244 = (CICC1851_resultStage_pixelStream_payload_245 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_245 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_246 = (CICC1851_resultStage_pixelStream_payload_247 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_247 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_248 = (CICC1851_resultStage_pixelStream_payload_249 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_249 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_when_SuperResolutionPart3_l1202 = (12'h003 + outRowCount_value);
  assign CICC1851_when_SuperResolutionPart3_l1205 = (12'h001 + outRowCount_value);
  assign CICC1851_when_SuperResolutionPart3_l1205_1 = (12'h002 + outPixelAddr_value);
  assign CICC1851_when_SuperResolutionPart3_l1205_2 = (12'h002 + outPixelAddr_value);
  assign CICC1851_when_SuperResolutionPart3_l1223 = {1'd0, outPixelAddr_value};
  assign CICC1851_when_SuperResolutionPart3_l1223_1 = (CICC1851_when_SuperResolutionPart3_l1223_2 - 13'h0002);
  assign CICC1851_when_SuperResolutionPart3_l1223_2 = (3'b100 * bmpWidth);
  assign CICC1851_when_SuperResolutionPart3_l1224 = {1'd0, outRowCount_value};
  assign CICC1851_when_SuperResolutionPart3_l1224_1 = (CICC1851_when_SuperResolutionPart3_l1224_2 - 13'h0002);
  assign CICC1851_when_SuperResolutionPart3_l1224_2 = (3'b100 * bmpHeight);
  assign CICC1851_lineBufferOne_port = passPixels_payload_pixel;
  assign CICC1851_lineBufferOne_port_1 = (passPixels_fire_6 && (bufferSwitch == 2'b00));
  assign CICC1851_lineBufferTwo_port = passPixels_payload_pixel;
  assign CICC1851_lineBufferTwo_port_1 = (passPixels_fire_7 && (bufferSwitch == 2'b01));
  assign CICC1851_lineBufferThree_port = passPixels_payload_pixel;
  assign CICC1851_lineBufferThree_port_1 = (passPixels_fire_8 && (bufferSwitch == 2'b10));
  assign CICC1851_validBufferOne_port = passPixels_payload_inpValid;
  assign CICC1851_validBufferOne_port_1 = (passPixels_fire_9 && (bufferSwitch == 2'b00));
  assign CICC1851_validBufferTwo_port = passPixels_payload_inpValid;
  assign CICC1851_validBufferTwo_port_1 = (passPixels_fire_10 && (bufferSwitch == 2'b01));
  assign CICC1851_validBufferThree_port = passPixels_payload_inpValid;
  assign CICC1851_validBufferThree_port_1 = (passPixels_fire_11 && (bufferSwitch == 2'b10));
  always @(posedge clk) begin
    if(CICC1851_lineBufferOne_port_1) begin
      lineBufferOne[bufferWAddr_value] <= CICC1851_lineBufferOne_port;
    end
  end

  always @(posedge clk) begin
    if(mainPixelAddrOneStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferOne_port1 <= lineBufferOne[mainPixelAddrOneStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(counterPixelAddrOneStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferOne_port2 <= lineBufferOne[counterPixelAddrOneStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(CICC1851_lineBufferTwo_port_1) begin
      lineBufferTwo[bufferWAddr_value] <= CICC1851_lineBufferTwo_port;
    end
  end

  always @(posedge clk) begin
    if(mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferTwo_port1 <= lineBufferTwo[mainPixelAddrTwoStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferTwo_port2 <= lineBufferTwo[counterPixelAddrTwoStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(CICC1851_lineBufferThree_port_1) begin
      lineBufferThree[bufferWAddr_value] <= CICC1851_lineBufferThree_port;
    end
  end

  always @(posedge clk) begin
    if(mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferThree_port1 <= lineBufferThree[mainPixelAddrThreeStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferThree_port2 <= lineBufferThree[counterPixelAddrThreeStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(CICC1851_validBufferOne_port_1) begin
      validBufferOne[bufferWAddr_value] <= CICC1851_validBufferOne_port;
    end
  end

  always @(posedge clk) begin
    if(mainValidAddrOneStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_validBufferOne_port1 <= validBufferOne[mainValidAddrOneStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(counterValidAddrOneStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_validBufferOne_port2 <= validBufferOne[counterValidAddrOneStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(CICC1851_validBufferTwo_port_1) begin
      validBufferTwo[bufferWAddr_value] <= CICC1851_validBufferTwo_port;
    end
  end

  always @(posedge clk) begin
    if(mainValidAddrTwoStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_validBufferTwo_port1 <= validBufferTwo[mainValidAddrTwoStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(counterValidAddrTwoStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_validBufferTwo_port2 <= validBufferTwo[counterValidAddrTwoStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(CICC1851_validBufferThree_port_1) begin
      validBufferThree[bufferWAddr_value] <= CICC1851_validBufferThree_port;
    end
  end

  always @(posedge clk) begin
    if(mainValidAddrThreeStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_validBufferThree_port1 <= validBufferThree[mainValidAddrThreeStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(counterValidAddrThreeStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_validBufferThree_port2 <= validBufferThree[counterValidAddrThreeStream_s2mPipe_m2sPipe_payload];
    end
  end

  StreamFork_3 diffStage_controlPipe_fork (
    .io_input_valid                                (diffStage_controlPipe_valid                                             ), //i
    .io_input_ready                                (diffStage_controlPipe_fork_io_input_ready                               ), //o
    .io_input_payload_frameStart                   (diffStage_controlPipe_payload_frameStart                                ), //i
    .io_input_payload_rowEnd                       (diffStage_controlPipe_payload_rowEnd                                    ), //i
    .io_input_payload_pipeValid                    (diffStage_controlPipe_payload_pipeValid                                 ), //i
    .io_input_payload_firstRow                     (diffStage_controlPipe_payload_firstRow                                  ), //i
    .io_input_payload_lastRow                      (diffStage_controlPipe_payload_lastRow                                   ), //i
    .io_input_payload_finalResult                  (diffStage_controlPipe_payload_finalResult                               ), //i
    .io_input_payload_mainCompare                  (diffStage_controlPipe_payload_mainCompare                               ), //i
    .io_input_payload_counterCompare               (diffStage_controlPipe_payload_counterCompare                            ), //i
    .io_input_payload_horizontalCompare            (diffStage_controlPipe_payload_horizontalCompare                         ), //i
    .io_input_payload_verticalCompare              (diffStage_controlPipe_payload_verticalCompare                           ), //i
    .io_input_payload_mainDiff                     (diffStage_controlPipe_payload_mainDiff[7:0]                             ), //i
    .io_input_payload_counterDiff                  (diffStage_controlPipe_payload_counterDiff[7:0]                          ), //i
    .io_input_payload_horizontalDiff               (diffStage_controlPipe_payload_horizontalDiff[7:0]                       ), //i
    .io_input_payload_verticalDiff                 (diffStage_controlPipe_payload_verticalDiff[7:0]                         ), //i
    .io_input_payload_isHorizontalMin              (diffStage_controlPipe_payload_isHorizontalMin                           ), //i
    .io_input_payload_minDiff                      (diffStage_controlPipe_payload_minDiff[7:0]                              ), //i
    .io_input_payload_currentPosition              (diffStage_controlPipe_payload_currentPosition[1:0]                      ), //i
    .io_input_payload_nextPosition                 (diffStage_controlPipe_payload_nextPosition[1:0]                         ), //i
    .io_input_payload_horizontalDirectionValid     (diffStage_controlPipe_payload_horizontalDirectionValid                  ), //i
    .io_input_payload_verticalDirectionValid       (diffStage_controlPipe_payload_verticalDirectionValid                    ), //i
    .io_input_payload_mainDirectionValid           (diffStage_controlPipe_payload_mainDirectionValid                        ), //i
    .io_input_payload_counterDirectionValid        (diffStage_controlPipe_payload_counterDirectionValid                     ), //i
    .io_input_payload_inValidMinDiff               (diffStage_controlPipe_payload_inValidMinDiff                            ), //i
    .io_outputs_0_valid                            (diffStage_controlPipe_fork_io_outputs_0_valid                           ), //o
    .io_outputs_0_ready                            (resultStage_controlPipeBeforePipe_ready                                 ), //i
    .io_outputs_0_payload_frameStart               (diffStage_controlPipe_fork_io_outputs_0_payload_frameStart              ), //o
    .io_outputs_0_payload_rowEnd                   (diffStage_controlPipe_fork_io_outputs_0_payload_rowEnd                  ), //o
    .io_outputs_0_payload_pipeValid                (diffStage_controlPipe_fork_io_outputs_0_payload_pipeValid               ), //o
    .io_outputs_0_payload_firstRow                 (diffStage_controlPipe_fork_io_outputs_0_payload_firstRow                ), //o
    .io_outputs_0_payload_lastRow                  (diffStage_controlPipe_fork_io_outputs_0_payload_lastRow                 ), //o
    .io_outputs_0_payload_finalResult              (diffStage_controlPipe_fork_io_outputs_0_payload_finalResult             ), //o
    .io_outputs_0_payload_mainCompare              (diffStage_controlPipe_fork_io_outputs_0_payload_mainCompare             ), //o
    .io_outputs_0_payload_counterCompare           (diffStage_controlPipe_fork_io_outputs_0_payload_counterCompare          ), //o
    .io_outputs_0_payload_horizontalCompare        (diffStage_controlPipe_fork_io_outputs_0_payload_horizontalCompare       ), //o
    .io_outputs_0_payload_verticalCompare          (diffStage_controlPipe_fork_io_outputs_0_payload_verticalCompare         ), //o
    .io_outputs_0_payload_mainDiff                 (diffStage_controlPipe_fork_io_outputs_0_payload_mainDiff[7:0]           ), //o
    .io_outputs_0_payload_counterDiff              (diffStage_controlPipe_fork_io_outputs_0_payload_counterDiff[7:0]        ), //o
    .io_outputs_0_payload_horizontalDiff           (diffStage_controlPipe_fork_io_outputs_0_payload_horizontalDiff[7:0]     ), //o
    .io_outputs_0_payload_verticalDiff             (diffStage_controlPipe_fork_io_outputs_0_payload_verticalDiff[7:0]       ), //o
    .io_outputs_0_payload_isHorizontalMin          (diffStage_controlPipe_fork_io_outputs_0_payload_isHorizontalMin         ), //o
    .io_outputs_0_payload_minDiff                  (diffStage_controlPipe_fork_io_outputs_0_payload_minDiff[7:0]            ), //o
    .io_outputs_0_payload_currentPosition          (diffStage_controlPipe_fork_io_outputs_0_payload_currentPosition[1:0]    ), //o
    .io_outputs_0_payload_nextPosition             (diffStage_controlPipe_fork_io_outputs_0_payload_nextPosition[1:0]       ), //o
    .io_outputs_0_payload_horizontalDirectionValid (diffStage_controlPipe_fork_io_outputs_0_payload_horizontalDirectionValid), //o
    .io_outputs_0_payload_verticalDirectionValid   (diffStage_controlPipe_fork_io_outputs_0_payload_verticalDirectionValid  ), //o
    .io_outputs_0_payload_mainDirectionValid       (diffStage_controlPipe_fork_io_outputs_0_payload_mainDirectionValid      ), //o
    .io_outputs_0_payload_counterDirectionValid    (diffStage_controlPipe_fork_io_outputs_0_payload_counterDirectionValid   ), //o
    .io_outputs_0_payload_inValidMinDiff           (diffStage_controlPipe_fork_io_outputs_0_payload_inValidMinDiff          ), //o
    .io_outputs_1_valid                            (diffStage_controlPipe_fork_io_outputs_1_valid                           ), //o
    .io_outputs_1_ready                            (resultStage_pixelStream_ready                                           ), //i
    .io_outputs_1_payload_frameStart               (diffStage_controlPipe_fork_io_outputs_1_payload_frameStart              ), //o
    .io_outputs_1_payload_rowEnd                   (diffStage_controlPipe_fork_io_outputs_1_payload_rowEnd                  ), //o
    .io_outputs_1_payload_pipeValid                (diffStage_controlPipe_fork_io_outputs_1_payload_pipeValid               ), //o
    .io_outputs_1_payload_firstRow                 (diffStage_controlPipe_fork_io_outputs_1_payload_firstRow                ), //o
    .io_outputs_1_payload_lastRow                  (diffStage_controlPipe_fork_io_outputs_1_payload_lastRow                 ), //o
    .io_outputs_1_payload_finalResult              (diffStage_controlPipe_fork_io_outputs_1_payload_finalResult             ), //o
    .io_outputs_1_payload_mainCompare              (diffStage_controlPipe_fork_io_outputs_1_payload_mainCompare             ), //o
    .io_outputs_1_payload_counterCompare           (diffStage_controlPipe_fork_io_outputs_1_payload_counterCompare          ), //o
    .io_outputs_1_payload_horizontalCompare        (diffStage_controlPipe_fork_io_outputs_1_payload_horizontalCompare       ), //o
    .io_outputs_1_payload_verticalCompare          (diffStage_controlPipe_fork_io_outputs_1_payload_verticalCompare         ), //o
    .io_outputs_1_payload_mainDiff                 (diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff[7:0]           ), //o
    .io_outputs_1_payload_counterDiff              (diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff[7:0]        ), //o
    .io_outputs_1_payload_horizontalDiff           (diffStage_controlPipe_fork_io_outputs_1_payload_horizontalDiff[7:0]     ), //o
    .io_outputs_1_payload_verticalDiff             (diffStage_controlPipe_fork_io_outputs_1_payload_verticalDiff[7:0]       ), //o
    .io_outputs_1_payload_isHorizontalMin          (diffStage_controlPipe_fork_io_outputs_1_payload_isHorizontalMin         ), //o
    .io_outputs_1_payload_minDiff                  (diffStage_controlPipe_fork_io_outputs_1_payload_minDiff[7:0]            ), //o
    .io_outputs_1_payload_currentPosition          (diffStage_controlPipe_fork_io_outputs_1_payload_currentPosition[1:0]    ), //o
    .io_outputs_1_payload_nextPosition             (diffStage_controlPipe_fork_io_outputs_1_payload_nextPosition[1:0]       ), //o
    .io_outputs_1_payload_horizontalDirectionValid (diffStage_controlPipe_fork_io_outputs_1_payload_horizontalDirectionValid), //o
    .io_outputs_1_payload_verticalDirectionValid   (diffStage_controlPipe_fork_io_outputs_1_payload_verticalDirectionValid  ), //o
    .io_outputs_1_payload_mainDirectionValid       (diffStage_controlPipe_fork_io_outputs_1_payload_mainDirectionValid      ), //o
    .io_outputs_1_payload_counterDirectionValid    (diffStage_controlPipe_fork_io_outputs_1_payload_counterDirectionValid   ), //o
    .io_outputs_1_payload_inValidMinDiff           (diffStage_controlPipe_fork_io_outputs_1_payload_inValidMinDiff          )  //o
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_8_BOOT : controlStateMachine_stateReg_string = "BOOT ";
      controlStateMachine_enumDef_8_HOLD : controlStateMachine_stateReg_string = "HOLD ";
      controlStateMachine_enumDef_8_PASS : controlStateMachine_stateReg_string = "PASS ";
      controlStateMachine_enumDef_8_EXTRA : controlStateMachine_stateReg_string = "EXTRA";
      default : controlStateMachine_stateReg_string = "?????";
    endcase
  end
  always @(*) begin
    case(controlStateMachine_stateNext)
      controlStateMachine_enumDef_8_BOOT : controlStateMachine_stateNext_string = "BOOT ";
      controlStateMachine_enumDef_8_HOLD : controlStateMachine_stateNext_string = "HOLD ";
      controlStateMachine_enumDef_8_PASS : controlStateMachine_stateNext_string = "PASS ";
      controlStateMachine_enumDef_8_EXTRA : controlStateMachine_stateNext_string = "EXTRA";
      default : controlStateMachine_stateNext_string = "?????";
    endcase
  end
  `endif

  always @(*) begin
    pixelsIn_ready = 1'b0;
    pixelsIn_ready = (! pixelsIn_rValid);
  end

  always @(*) begin
    pixelsOut_valid = 1'b0;
    pixelsOut_valid = pixelsStream_s2mPipe_m2sPipe_valid;
  end

  always @(*) begin
    pixelsOut_payload_pixel = 8'h0;
    pixelsOut_payload_pixel = pixelsStream_s2mPipe_m2sPipe_payload_pixel;
  end

  always @(*) begin
    pixelsOut_payload_frameStart = 1'b0;
    pixelsOut_payload_frameStart = pixelsStream_s2mPipe_m2sPipe_payload_frameStart;
  end

  always @(*) begin
    pixelsOut_payload_rowEnd = 1'b0;
    pixelsOut_payload_rowEnd = pixelsStream_s2mPipe_m2sPipe_payload_rowEnd;
  end

  always @(*) begin
    inpThreeDoneOut = 1'b0;
    inpThreeDoneOut = inpThreeDone;
  end

  assign when_SuperResolutionPart3_l72 = (startIn && (! startIn_regNext));
  assign when_SuperResolutionPart3_l75 = (! startIn);
  assign when_SuperResolutionPart3_l78 = (startIn && (! readDone));
  assign when_SuperResolutionPart3_l78_1 = (! startIn);
  assign when_SuperResolutionPart3_l93 = (! startIn);
  assign when_SuperResolutionPart3_l96 = (! startIn);
  always @(*) begin
    bufferRowCount_willIncrement = 1'b0;
    if(when_SuperResolutionPart3_l230) begin
      if(!bufferReachFinalRow) begin
        bufferRowCount_willIncrement = 1'b1;
      end
    end
  end

  always @(*) begin
    bufferRowCount_willClear = 1'b0;
    if(when_SuperResolutionPart3_l230) begin
      if(bufferReachFinalRow) begin
        bufferRowCount_willClear = 1'b1;
      end
    end
  end

  assign bufferRowCount_willOverflowIfInc = (bufferRowCount_value == 12'h870);
  assign bufferRowCount_willOverflow = (bufferRowCount_willOverflowIfInc && bufferRowCount_willIncrement);
  always @(*) begin
    if(bufferRowCount_willOverflow) begin
      bufferRowCount_valueNext = 12'h0;
    end else begin
      bufferRowCount_valueNext = (bufferRowCount_value + CICC1851_bufferRowCount_valueNext);
    end
    if(bufferRowCount_willClear) begin
      bufferRowCount_valueNext = 12'h0;
    end
  end

  assign when_SuperResolutionPart3_l102 = ((startIn && (! holdBuffer)) && (! writeDone));
  assign when_SuperResolutionPart3_l102_1 = (((! startIn) || holdBuffer) || writeDone);
  always @(*) begin
    bufferWAddr_willIncrement = 1'b0;
    if(passPixels_fire_12) begin
      if(!passPixels_payload_rowEnd) begin
        bufferWAddr_willIncrement = 1'b1;
      end
    end
  end

  always @(*) begin
    bufferWAddr_willClear = 1'b0;
    if(passPixels_fire_12) begin
      if(passPixels_payload_rowEnd) begin
        bufferWAddr_willClear = 1'b1;
      end
    end
  end

  assign bufferWAddr_willOverflowIfInc = (bufferWAddr_value == 12'heff);
  assign bufferWAddr_willOverflow = (bufferWAddr_willOverflowIfInc && bufferWAddr_willIncrement);
  always @(*) begin
    if(bufferWAddr_willOverflow) begin
      bufferWAddr_valueNext = 12'h0;
    end else begin
      bufferWAddr_valueNext = (bufferWAddr_value + CICC1851_bufferWAddr_valueNext);
    end
    if(bufferWAddr_willClear) begin
      bufferWAddr_valueNext = 12'h0;
    end
  end

  always @(*) begin
    outPixelAddr_willIncrement = 1'b0;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_8_HOLD : begin
      end
      controlStateMachine_enumDef_8_PASS : begin
      end
      controlStateMachine_enumDef_8_EXTRA : begin
        if(controlStream_fire_6) begin
          if(!outReachRowEnd) begin
            outPixelAddr_willIncrement = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outPixelAddr_willClear = 1'b0;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_8_HOLD : begin
      end
      controlStateMachine_enumDef_8_PASS : begin
      end
      controlStateMachine_enumDef_8_EXTRA : begin
        if(controlStream_fire_6) begin
          if(outReachRowEnd) begin
            outPixelAddr_willClear = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign outPixelAddr_willOverflowIfInc = (outPixelAddr_value == 12'heff);
  assign outPixelAddr_willOverflow = (outPixelAddr_willOverflowIfInc && outPixelAddr_willIncrement);
  always @(*) begin
    if(outPixelAddr_willOverflow) begin
      outPixelAddr_valueNext = 12'h0;
    end else begin
      outPixelAddr_valueNext = (outPixelAddr_value + CICC1851_outPixelAddr_valueNext);
    end
    if(outPixelAddr_willClear) begin
      outPixelAddr_valueNext = 12'h0;
    end
  end

  always @(*) begin
    outRowCount_willIncrement = 1'b0;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_8_HOLD : begin
      end
      controlStateMachine_enumDef_8_PASS : begin
      end
      controlStateMachine_enumDef_8_EXTRA : begin
        if(when_SuperResolutionPart3_l1226) begin
          if(!outReachFinalRow) begin
            outRowCount_willIncrement = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outRowCount_willClear = 1'b0;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_8_HOLD : begin
      end
      controlStateMachine_enumDef_8_PASS : begin
      end
      controlStateMachine_enumDef_8_EXTRA : begin
        if(when_SuperResolutionPart3_l1226) begin
          if(outReachFinalRow) begin
            outRowCount_willClear = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign outRowCount_willOverflowIfInc = (outRowCount_value == 12'h870);
  assign outRowCount_willOverflow = (outRowCount_willOverflowIfInc && outRowCount_willIncrement);
  always @(*) begin
    if(outRowCount_willOverflow) begin
      outRowCount_valueNext = 12'h0;
    end else begin
      outRowCount_valueNext = (outRowCount_value + CICC1851_outRowCount_valueNext);
    end
    if(outRowCount_willClear) begin
      outRowCount_valueNext = 12'h0;
    end
  end

  always @(*) begin
    alreadySendRow_willIncrement = 1'b0;
    if(pixelsOut_fire_2) begin
      if(alreadyReachRowEnd) begin
        if(!alreadyReachFinalRow) begin
          alreadySendRow_willIncrement = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    alreadySendRow_willClear = 1'b0;
    if(pixelsOut_fire_2) begin
      if(alreadyReachRowEnd) begin
        if(alreadyReachFinalRow) begin
          alreadySendRow_willClear = 1'b1;
        end
      end
    end
  end

  assign alreadySendRow_willOverflowIfInc = (alreadySendRow_value == 12'h870);
  assign alreadySendRow_willOverflow = (alreadySendRow_willOverflowIfInc && alreadySendRow_willIncrement);
  always @(*) begin
    if(alreadySendRow_willOverflow) begin
      alreadySendRow_valueNext = 12'h0;
    end else begin
      alreadySendRow_valueNext = (alreadySendRow_value + CICC1851_alreadySendRow_valueNext);
    end
    if(alreadySendRow_willClear) begin
      alreadySendRow_valueNext = 12'h0;
    end
  end

  always @(*) begin
    alreadySendCountInRow_willIncrement = 1'b0;
    if(pixelsOut_fire_2) begin
      if(!alreadyReachRowEnd) begin
        alreadySendCountInRow_willIncrement = 1'b1;
      end
    end
  end

  always @(*) begin
    alreadySendCountInRow_willClear = 1'b0;
    if(pixelsOut_fire_2) begin
      if(alreadyReachRowEnd) begin
        alreadySendCountInRow_willClear = 1'b1;
      end
    end
  end

  assign alreadySendCountInRow_willOverflowIfInc = (alreadySendCountInRow_value == 12'heff);
  assign alreadySendCountInRow_willOverflow = (alreadySendCountInRow_willOverflowIfInc && alreadySendCountInRow_willIncrement);
  always @(*) begin
    if(alreadySendCountInRow_willOverflow) begin
      alreadySendCountInRow_valueNext = 12'h0;
    end else begin
      alreadySendCountInRow_valueNext = (alreadySendCountInRow_value + CICC1851_alreadySendCountInRow_valueNext);
    end
    if(alreadySendCountInRow_willClear) begin
      alreadySendCountInRow_valueNext = 12'h0;
    end
  end

  assign when_SuperResolutionPart3_l154 = ((! startRead) || ((! startIn) && startIn_regNext_1));
  always @(*) begin
    mainAddrOne = outPixelAddr_value;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_8_HOLD : begin
      end
      controlStateMachine_enumDef_8_PASS : begin
        if(when_SuperResolutionPart3_l1168) begin
          mainAddrOne = (12'h001 + outPixelAddr_value);
        end else begin
          mainAddrOne = (outPixelAddr_value - 12'h001);
        end
      end
      controlStateMachine_enumDef_8_EXTRA : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    counterAddrOne = outPixelAddr_value;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_8_HOLD : begin
      end
      controlStateMachine_enumDef_8_PASS : begin
        if(outReachRowEnd) begin
          counterAddrOne = (outPixelAddr_value - 12'h001);
        end else begin
          counterAddrOne = (12'h001 + outPixelAddr_value);
        end
      end
      controlStateMachine_enumDef_8_EXTRA : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    mainAddrTwo = outPixelAddr_value;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_8_HOLD : begin
      end
      controlStateMachine_enumDef_8_PASS : begin
        if(when_SuperResolutionPart3_l1168) begin
          mainAddrTwo = (12'h001 + outPixelAddr_value);
        end else begin
          mainAddrTwo = (outPixelAddr_value - 12'h001);
        end
      end
      controlStateMachine_enumDef_8_EXTRA : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    counterAddrTwo = outPixelAddr_value;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_8_HOLD : begin
      end
      controlStateMachine_enumDef_8_PASS : begin
        if(outReachRowEnd) begin
          counterAddrTwo = (outPixelAddr_value - 12'h001);
        end else begin
          counterAddrTwo = (12'h001 + outPixelAddr_value);
        end
      end
      controlStateMachine_enumDef_8_EXTRA : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    mainAddrThree = outPixelAddr_value;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_8_HOLD : begin
      end
      controlStateMachine_enumDef_8_PASS : begin
        if(when_SuperResolutionPart3_l1168) begin
          mainAddrThree = (12'h001 + outPixelAddr_value);
        end else begin
          mainAddrThree = (outPixelAddr_value - 12'h001);
        end
      end
      controlStateMachine_enumDef_8_EXTRA : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    counterAddrThree = outPixelAddr_value;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_8_HOLD : begin
      end
      controlStateMachine_enumDef_8_PASS : begin
        if(outReachRowEnd) begin
          counterAddrThree = (outPixelAddr_value - 12'h001);
        end else begin
          counterAddrThree = (12'h001 + outPixelAddr_value);
        end
      end
      controlStateMachine_enumDef_8_EXTRA : begin
      end
      default : begin
      end
    endcase
  end

  assign validStream_valid = 1'b1;
  assign CICC1851_controls_frameStart = 60'h0;
  always @(*) begin
    controls_frameStart = CICC1851_controls_frameStart[0];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_8_HOLD : begin
      end
      controlStateMachine_enumDef_8_PASS : begin
        if(frameStart) begin
          controls_frameStart = 1'b1;
        end
      end
      controlStateMachine_enumDef_8_EXTRA : begin
        if(frameStart) begin
          controls_frameStart = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_rowEnd = CICC1851_controls_frameStart[1];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_8_HOLD : begin
      end
      controlStateMachine_enumDef_8_PASS : begin
        if(outReachRowEnd) begin
          controls_rowEnd = 1'b1;
        end
      end
      controlStateMachine_enumDef_8_EXTRA : begin
        if(outReachRowEnd) begin
          controls_rowEnd = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_pipeValid = CICC1851_controls_frameStart[2];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_8_HOLD : begin
      end
      controlStateMachine_enumDef_8_PASS : begin
        controls_pipeValid = 1'b1;
      end
      controlStateMachine_enumDef_8_EXTRA : begin
        controls_pipeValid = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_firstRow = CICC1851_controls_frameStart[3];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_8_HOLD : begin
      end
      controlStateMachine_enumDef_8_PASS : begin
        if(when_SuperResolutionPart3_l1188) begin
          controls_firstRow = 1'b1;
        end
      end
      controlStateMachine_enumDef_8_EXTRA : begin
        if(when_SuperResolutionPart3_l1217) begin
          controls_firstRow = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_lastRow = CICC1851_controls_frameStart[4];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_8_HOLD : begin
      end
      controlStateMachine_enumDef_8_PASS : begin
        if(outReachFinalRow) begin
          controls_lastRow = 1'b1;
        end
      end
      controlStateMachine_enumDef_8_EXTRA : begin
        if(outReachFinalRow) begin
          controls_lastRow = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_finalResult = CICC1851_controls_frameStart[5];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_8_HOLD : begin
      end
      controlStateMachine_enumDef_8_PASS : begin
      end
      controlStateMachine_enumDef_8_EXTRA : begin
        controls_finalResult = 1'b1;
      end
      default : begin
      end
    endcase
  end

  assign controls_mainCompare = CICC1851_controls_frameStart[6];
  assign controls_counterCompare = CICC1851_controls_frameStart[7];
  assign controls_horizontalCompare = CICC1851_controls_frameStart[8];
  assign controls_verticalCompare = CICC1851_controls_frameStart[9];
  assign controls_mainDiff = CICC1851_controls_frameStart[17 : 10];
  assign controls_counterDiff = CICC1851_controls_frameStart[25 : 18];
  assign controls_horizontalDiff = CICC1851_controls_frameStart[33 : 26];
  assign controls_verticalDiff = CICC1851_controls_frameStart[41 : 34];
  assign controls_isHorizontalMin = CICC1851_controls_frameStart[42];
  assign controls_minDiff = CICC1851_controls_frameStart[50 : 43];
  always @(*) begin
    controls_currentPosition = CICC1851_controls_frameStart[52 : 51];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_8_HOLD : begin
      end
      controlStateMachine_enumDef_8_PASS : begin
        controls_currentPosition = currentRowBuffer;
      end
      controlStateMachine_enumDef_8_EXTRA : begin
        controls_currentPosition = currentRowBuffer;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_nextPosition = CICC1851_controls_frameStart[54 : 53];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_8_HOLD : begin
      end
      controlStateMachine_enumDef_8_PASS : begin
        controls_nextPosition = nextRowBuffer;
      end
      controlStateMachine_enumDef_8_EXTRA : begin
        controls_nextPosition = nextRowBuffer;
      end
      default : begin
      end
    endcase
  end

  assign controls_horizontalDirectionValid = CICC1851_controls_frameStart[55];
  assign controls_verticalDirectionValid = CICC1851_controls_frameStart[56];
  assign controls_mainDirectionValid = CICC1851_controls_frameStart[57];
  assign controls_counterDirectionValid = CICC1851_controls_frameStart[58];
  assign controls_inValidMinDiff = CICC1851_controls_frameStart[59];
  always @(*) begin
    validStream_ready = (controlStream_ready && startRead);
    validStream_ready = (mainPixelAddrOneStream_ready && startRead);
    validStream_ready = (counterPixelAddrOneStream_ready && startRead);
    validStream_ready = (mainPixelAddrTwoStream_ready && startRead);
    validStream_ready = (counterPixelAddrTwoStream_ready && startRead);
    validStream_ready = (mainPixelAddrThreeStream_ready && startRead);
    validStream_ready = (counterPixelAddrThreeStream_ready && startRead);
    validStream_ready = (mainValidAddrOneStream_ready && startRead);
    validStream_ready = (counterValidAddrOneStream_ready && startRead);
    validStream_ready = (mainValidAddrTwoStream_ready && startRead);
    validStream_ready = (counterValidAddrTwoStream_ready && startRead);
    validStream_ready = (mainValidAddrThreeStream_ready && startRead);
    validStream_ready = (counterValidAddrThreeStream_ready && startRead);
  end

  assign controlStream_valid = (validStream_valid && startRead);
  assign controlStream_payload_frameStart = controls_frameStart;
  assign controlStream_payload_rowEnd = controls_rowEnd;
  assign controlStream_payload_pipeValid = controls_pipeValid;
  assign controlStream_payload_firstRow = controls_firstRow;
  assign controlStream_payload_lastRow = controls_lastRow;
  assign controlStream_payload_finalResult = controls_finalResult;
  assign controlStream_payload_mainCompare = controls_mainCompare;
  assign controlStream_payload_counterCompare = controls_counterCompare;
  assign controlStream_payload_horizontalCompare = controls_horizontalCompare;
  assign controlStream_payload_verticalCompare = controls_verticalCompare;
  assign controlStream_payload_mainDiff = controls_mainDiff;
  assign controlStream_payload_counterDiff = controls_counterDiff;
  assign controlStream_payload_horizontalDiff = controls_horizontalDiff;
  assign controlStream_payload_verticalDiff = controls_verticalDiff;
  assign controlStream_payload_isHorizontalMin = controls_isHorizontalMin;
  assign controlStream_payload_minDiff = controls_minDiff;
  assign controlStream_payload_currentPosition = controls_currentPosition;
  assign controlStream_payload_nextPosition = controls_nextPosition;
  assign controlStream_payload_horizontalDirectionValid = controls_horizontalDirectionValid;
  assign controlStream_payload_verticalDirectionValid = controls_verticalDirectionValid;
  assign controlStream_payload_mainDirectionValid = controls_mainDirectionValid;
  assign controlStream_payload_counterDirectionValid = controls_counterDirectionValid;
  assign controlStream_payload_inValidMinDiff = controls_inValidMinDiff;
  assign mainPixelAddrOneStream_valid = (validStream_valid && startRead);
  assign mainPixelAddrOneStream_payload = mainAddrOne;
  assign counterPixelAddrOneStream_valid = (validStream_valid && startRead);
  assign counterPixelAddrOneStream_payload = counterAddrOne;
  assign mainPixelAddrTwoStream_valid = (validStream_valid && startRead);
  assign mainPixelAddrTwoStream_payload = mainAddrTwo;
  assign counterPixelAddrTwoStream_valid = (validStream_valid && startRead);
  assign counterPixelAddrTwoStream_payload = counterAddrTwo;
  assign mainPixelAddrThreeStream_valid = (validStream_valid && startRead);
  assign mainPixelAddrThreeStream_payload = mainAddrThree;
  assign counterPixelAddrThreeStream_valid = (validStream_valid && startRead);
  assign counterPixelAddrThreeStream_payload = counterAddrThree;
  assign mainValidAddrOneStream_valid = (validStream_valid && startRead);
  assign mainValidAddrOneStream_payload = mainAddrOne;
  assign counterValidAddrOneStream_valid = (validStream_valid && startRead);
  assign counterValidAddrOneStream_payload = counterAddrOne;
  assign mainValidAddrTwoStream_valid = (validStream_valid && startRead);
  assign mainValidAddrTwoStream_payload = mainAddrTwo;
  assign counterValidAddrTwoStream_valid = (validStream_valid && startRead);
  assign counterValidAddrTwoStream_payload = counterAddrTwo;
  assign mainValidAddrThreeStream_valid = (validStream_valid && startRead);
  assign mainValidAddrThreeStream_payload = mainAddrThree;
  assign counterValidAddrThreeStream_valid = (validStream_valid && startRead);
  assign counterValidAddrThreeStream_payload = counterAddrThree;
  assign pixelsIn_s2mPipe_valid = (pixelsIn_valid || pixelsIn_rValid);
  assign pixelsIn_s2mPipe_payload_pixel = (pixelsIn_rValid ? pixelsIn_rData_pixel : pixelsIn_payload_pixel);
  assign pixelsIn_s2mPipe_payload_frameStart = (pixelsIn_rValid ? pixelsIn_rData_frameStart : pixelsIn_payload_frameStart);
  assign pixelsIn_s2mPipe_payload_rowEnd = (pixelsIn_rValid ? pixelsIn_rData_rowEnd : pixelsIn_payload_rowEnd);
  assign pixelsIn_s2mPipe_payload_inpValid = (pixelsIn_rValid ? pixelsIn_rData_inpValid : pixelsIn_payload_inpValid);
  always @(*) begin
    pixelsIn_s2mPipe_ready = pixelsIn_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368) begin
      pixelsIn_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368 = (! pixelsIn_s2mPipe_m2sPipe_valid);
  assign pixelsIn_s2mPipe_m2sPipe_valid = pixelsIn_s2mPipe_rValid;
  assign pixelsIn_s2mPipe_m2sPipe_payload_pixel = pixelsIn_s2mPipe_rData_pixel;
  assign pixelsIn_s2mPipe_m2sPipe_payload_frameStart = pixelsIn_s2mPipe_rData_frameStart;
  assign pixelsIn_s2mPipe_m2sPipe_payload_rowEnd = pixelsIn_s2mPipe_rData_rowEnd;
  assign pixelsIn_s2mPipe_m2sPipe_payload_inpValid = pixelsIn_s2mPipe_rData_inpValid;
  assign passPixels_valid = (pixelsIn_s2mPipe_m2sPipe_valid && bufferEnable);
  assign pixelsIn_s2mPipe_m2sPipe_ready = (passPixels_ready && bufferEnable);
  assign passPixels_payload_pixel = pixelsIn_s2mPipe_m2sPipe_payload_pixel;
  assign passPixels_payload_frameStart = pixelsIn_s2mPipe_m2sPipe_payload_frameStart;
  assign passPixels_payload_rowEnd = pixelsIn_s2mPipe_m2sPipe_payload_rowEnd;
  assign passPixels_payload_inpValid = pixelsIn_s2mPipe_m2sPipe_payload_inpValid;
  assign passPixels_ready = 1'b1;
  assign passPixels_fire = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart3_l226 = ((CICC1851_when_SuperResolutionPart3_l226 == CICC1851_when_SuperResolutionPart3_l226_1) && passPixels_fire);
  assign passPixels_fire_1 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart3_l227 = (((CICC1851_when_SuperResolutionPart3_l227 == CICC1851_when_SuperResolutionPart3_l227_1) && bufferReachRowEnd) && passPixels_fire_1);
  assign passPixels_fire_2 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart3_l230 = (passPixels_payload_rowEnd && passPixels_fire_2);
  assign passPixels_fire_3 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart3_l243 = (passPixels_payload_rowEnd && passPixels_fire_3);
  assign when_SuperResolutionPart3_l244 = (bufferSwitch == 2'b10);
  assign passPixels_fire_4 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart3_l251 = (((12'h002 <= bufferRowCount_value) && passPixels_payload_rowEnd) && passPixels_fire_4);
  assign when_SuperResolutionPart3_l255 = (bufferReachFinalRow && bufferReachRowEnd);
  assign passPixels_fire_5 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart3_l262 = (passPixels_payload_frameStart && passPixels_fire_5);
  assign pixelsOut_fire = (pixelsOut_valid && pixelsOut_ready);
  assign when_SuperResolutionPart3_l270 = ((CICC1851_when_SuperResolutionPart3_l270 == CICC1851_when_SuperResolutionPart3_l270_1) && pixelsOut_fire);
  assign pixelsOut_fire_1 = (pixelsOut_valid && pixelsOut_ready);
  assign when_SuperResolutionPart3_l271 = (((CICC1851_when_SuperResolutionPart3_l271 == CICC1851_when_SuperResolutionPart3_l271_1) && alreadyReachRowEnd) && pixelsOut_fire_1);
  assign pixelsOut_fire_2 = (pixelsOut_valid && pixelsOut_ready);
  assign pixelsOut_fire_3 = (pixelsOut_valid && pixelsOut_ready);
  assign when_SuperResolutionPart3_l282 = ((alreadyReachFinalRow && alreadyReachRowEnd) && pixelsOut_fire_3);
  assign passPixels_fire_6 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_7 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_8 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_9 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_10 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_11 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_12 = (passPixels_valid && passPixels_ready);
  assign mainPixelAddrOneStream_ready = (! mainPixelAddrOneStream_rValid);
  assign mainPixelAddrOneStream_s2mPipe_valid = (mainPixelAddrOneStream_valid || mainPixelAddrOneStream_rValid);
  assign mainPixelAddrOneStream_s2mPipe_payload = (mainPixelAddrOneStream_rValid ? mainPixelAddrOneStream_rData : mainPixelAddrOneStream_payload);
  always @(*) begin
    mainPixelAddrOneStream_s2mPipe_ready = mainPixelAddrOneStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_1) begin
      mainPixelAddrOneStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_1 = (! mainPixelAddrOneStream_s2mPipe_m2sPipe_valid);
  assign mainPixelAddrOneStream_s2mPipe_m2sPipe_valid = mainPixelAddrOneStream_s2mPipe_rValid;
  assign mainPixelAddrOneStream_s2mPipe_m2sPipe_payload = mainPixelAddrOneStream_s2mPipe_rData;
  assign mainPixelAddrOneStream_s2mPipe_m2sPipe_ready = ((! CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready) || CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready = CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_mainOnePixelStream_payload = CICC1851_lineBufferOne_port1;
  assign CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_1 = readStage_mainOnePixelStream_ready;
    if(when_Stream_l368_2) begin
      CICC1851_1 = 1'b1;
    end
  end

  assign when_Stream_l368_2 = (! readStage_mainOnePixelStream_valid);
  assign readStage_mainOnePixelStream_valid = CICC1851_readStage_mainOnePixelStream_valid;
  assign readStage_mainOnePixelStream_payload = CICC1851_readStage_mainOnePixelStream_payload_2;
  assign counterPixelAddrOneStream_ready = (! counterPixelAddrOneStream_rValid);
  assign counterPixelAddrOneStream_s2mPipe_valid = (counterPixelAddrOneStream_valid || counterPixelAddrOneStream_rValid);
  assign counterPixelAddrOneStream_s2mPipe_payload = (counterPixelAddrOneStream_rValid ? counterPixelAddrOneStream_rData : counterPixelAddrOneStream_payload);
  always @(*) begin
    counterPixelAddrOneStream_s2mPipe_ready = counterPixelAddrOneStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_3) begin
      counterPixelAddrOneStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_3 = (! counterPixelAddrOneStream_s2mPipe_m2sPipe_valid);
  assign counterPixelAddrOneStream_s2mPipe_m2sPipe_valid = counterPixelAddrOneStream_s2mPipe_rValid;
  assign counterPixelAddrOneStream_s2mPipe_m2sPipe_payload = counterPixelAddrOneStream_s2mPipe_rData;
  assign counterPixelAddrOneStream_s2mPipe_m2sPipe_ready = ((! CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready) || CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready = CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_counterOnePixelStream_payload = CICC1851_lineBufferOne_port2;
  assign CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_2 = readStage_counterOnePixelStream_ready;
    if(when_Stream_l368_4) begin
      CICC1851_2 = 1'b1;
    end
  end

  assign when_Stream_l368_4 = (! readStage_counterOnePixelStream_valid);
  assign readStage_counterOnePixelStream_valid = CICC1851_readStage_counterOnePixelStream_valid;
  assign readStage_counterOnePixelStream_payload = CICC1851_readStage_counterOnePixelStream_payload_2;
  assign mainPixelAddrTwoStream_ready = (! mainPixelAddrTwoStream_rValid);
  assign mainPixelAddrTwoStream_s2mPipe_valid = (mainPixelAddrTwoStream_valid || mainPixelAddrTwoStream_rValid);
  assign mainPixelAddrTwoStream_s2mPipe_payload = (mainPixelAddrTwoStream_rValid ? mainPixelAddrTwoStream_rData : mainPixelAddrTwoStream_payload);
  always @(*) begin
    mainPixelAddrTwoStream_s2mPipe_ready = mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_5) begin
      mainPixelAddrTwoStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_5 = (! mainPixelAddrTwoStream_s2mPipe_m2sPipe_valid);
  assign mainPixelAddrTwoStream_s2mPipe_m2sPipe_valid = mainPixelAddrTwoStream_s2mPipe_rValid;
  assign mainPixelAddrTwoStream_s2mPipe_m2sPipe_payload = mainPixelAddrTwoStream_s2mPipe_rData;
  assign mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready = ((! CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready) || CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready = CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_mainTwoPixelStream_payload = CICC1851_lineBufferTwo_port1;
  assign CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_3 = readStage_mainTwoPixelStream_ready;
    if(when_Stream_l368_6) begin
      CICC1851_3 = 1'b1;
    end
  end

  assign when_Stream_l368_6 = (! readStage_mainTwoPixelStream_valid);
  assign readStage_mainTwoPixelStream_valid = CICC1851_readStage_mainTwoPixelStream_valid;
  assign readStage_mainTwoPixelStream_payload = CICC1851_readStage_mainTwoPixelStream_payload_2;
  assign counterPixelAddrTwoStream_ready = (! counterPixelAddrTwoStream_rValid);
  assign counterPixelAddrTwoStream_s2mPipe_valid = (counterPixelAddrTwoStream_valid || counterPixelAddrTwoStream_rValid);
  assign counterPixelAddrTwoStream_s2mPipe_payload = (counterPixelAddrTwoStream_rValid ? counterPixelAddrTwoStream_rData : counterPixelAddrTwoStream_payload);
  always @(*) begin
    counterPixelAddrTwoStream_s2mPipe_ready = counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_7) begin
      counterPixelAddrTwoStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_7 = (! counterPixelAddrTwoStream_s2mPipe_m2sPipe_valid);
  assign counterPixelAddrTwoStream_s2mPipe_m2sPipe_valid = counterPixelAddrTwoStream_s2mPipe_rValid;
  assign counterPixelAddrTwoStream_s2mPipe_m2sPipe_payload = counterPixelAddrTwoStream_s2mPipe_rData;
  assign counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready = ((! CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready) || CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready = CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_counterTwoPixelStream_payload = CICC1851_lineBufferTwo_port2;
  assign CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_4 = readStage_counterTwoPixelStream_ready;
    if(when_Stream_l368_8) begin
      CICC1851_4 = 1'b1;
    end
  end

  assign when_Stream_l368_8 = (! readStage_counterTwoPixelStream_valid);
  assign readStage_counterTwoPixelStream_valid = CICC1851_readStage_counterTwoPixelStream_valid;
  assign readStage_counterTwoPixelStream_payload = CICC1851_readStage_counterTwoPixelStream_payload_2;
  assign mainPixelAddrThreeStream_ready = (! mainPixelAddrThreeStream_rValid);
  assign mainPixelAddrThreeStream_s2mPipe_valid = (mainPixelAddrThreeStream_valid || mainPixelAddrThreeStream_rValid);
  assign mainPixelAddrThreeStream_s2mPipe_payload = (mainPixelAddrThreeStream_rValid ? mainPixelAddrThreeStream_rData : mainPixelAddrThreeStream_payload);
  always @(*) begin
    mainPixelAddrThreeStream_s2mPipe_ready = mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_9) begin
      mainPixelAddrThreeStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_9 = (! mainPixelAddrThreeStream_s2mPipe_m2sPipe_valid);
  assign mainPixelAddrThreeStream_s2mPipe_m2sPipe_valid = mainPixelAddrThreeStream_s2mPipe_rValid;
  assign mainPixelAddrThreeStream_s2mPipe_m2sPipe_payload = mainPixelAddrThreeStream_s2mPipe_rData;
  assign mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready = ((! CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready) || CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready = CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_mainThreePixelStream_payload = CICC1851_lineBufferThree_port1;
  assign CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_5 = readStage_mainThreePixelStream_ready;
    if(when_Stream_l368_10) begin
      CICC1851_5 = 1'b1;
    end
  end

  assign when_Stream_l368_10 = (! readStage_mainThreePixelStream_valid);
  assign readStage_mainThreePixelStream_valid = CICC1851_readStage_mainThreePixelStream_valid;
  assign readStage_mainThreePixelStream_payload = CICC1851_readStage_mainThreePixelStream_payload_2;
  assign counterPixelAddrThreeStream_ready = (! counterPixelAddrThreeStream_rValid);
  assign counterPixelAddrThreeStream_s2mPipe_valid = (counterPixelAddrThreeStream_valid || counterPixelAddrThreeStream_rValid);
  assign counterPixelAddrThreeStream_s2mPipe_payload = (counterPixelAddrThreeStream_rValid ? counterPixelAddrThreeStream_rData : counterPixelAddrThreeStream_payload);
  always @(*) begin
    counterPixelAddrThreeStream_s2mPipe_ready = counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_11) begin
      counterPixelAddrThreeStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_11 = (! counterPixelAddrThreeStream_s2mPipe_m2sPipe_valid);
  assign counterPixelAddrThreeStream_s2mPipe_m2sPipe_valid = counterPixelAddrThreeStream_s2mPipe_rValid;
  assign counterPixelAddrThreeStream_s2mPipe_m2sPipe_payload = counterPixelAddrThreeStream_s2mPipe_rData;
  assign counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready = ((! CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready) || CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready = CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_counterThreePixelStream_payload = CICC1851_lineBufferThree_port2;
  assign CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_6 = readStage_counterThreePixelStream_ready;
    if(when_Stream_l368_12) begin
      CICC1851_6 = 1'b1;
    end
  end

  assign when_Stream_l368_12 = (! readStage_counterThreePixelStream_valid);
  assign readStage_counterThreePixelStream_valid = CICC1851_readStage_counterThreePixelStream_valid;
  assign readStage_counterThreePixelStream_payload = CICC1851_readStage_counterThreePixelStream_payload_2;
  assign mainValidAddrOneStream_ready = (! mainValidAddrOneStream_rValid);
  assign mainValidAddrOneStream_s2mPipe_valid = (mainValidAddrOneStream_valid || mainValidAddrOneStream_rValid);
  assign mainValidAddrOneStream_s2mPipe_payload = (mainValidAddrOneStream_rValid ? mainValidAddrOneStream_rData : mainValidAddrOneStream_payload);
  always @(*) begin
    mainValidAddrOneStream_s2mPipe_ready = mainValidAddrOneStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_13) begin
      mainValidAddrOneStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_13 = (! mainValidAddrOneStream_s2mPipe_m2sPipe_valid);
  assign mainValidAddrOneStream_s2mPipe_m2sPipe_valid = mainValidAddrOneStream_s2mPipe_rValid;
  assign mainValidAddrOneStream_s2mPipe_m2sPipe_payload = mainValidAddrOneStream_s2mPipe_rData;
  assign mainValidAddrOneStream_s2mPipe_m2sPipe_ready = ((! CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready) || CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready = CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_mainOneValidStream_payload = CICC1851_validBufferOne_port1[0];
  assign CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_7 = readStage_mainOneValidStream_ready;
    if(when_Stream_l368_14) begin
      CICC1851_7 = 1'b1;
    end
  end

  assign when_Stream_l368_14 = (! readStage_mainOneValidStream_valid);
  assign readStage_mainOneValidStream_valid = CICC1851_readStage_mainOneValidStream_valid;
  assign readStage_mainOneValidStream_payload = CICC1851_readStage_mainOneValidStream_payload_2;
  assign counterValidAddrOneStream_ready = (! counterValidAddrOneStream_rValid);
  assign counterValidAddrOneStream_s2mPipe_valid = (counterValidAddrOneStream_valid || counterValidAddrOneStream_rValid);
  assign counterValidAddrOneStream_s2mPipe_payload = (counterValidAddrOneStream_rValid ? counterValidAddrOneStream_rData : counterValidAddrOneStream_payload);
  always @(*) begin
    counterValidAddrOneStream_s2mPipe_ready = counterValidAddrOneStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_15) begin
      counterValidAddrOneStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_15 = (! counterValidAddrOneStream_s2mPipe_m2sPipe_valid);
  assign counterValidAddrOneStream_s2mPipe_m2sPipe_valid = counterValidAddrOneStream_s2mPipe_rValid;
  assign counterValidAddrOneStream_s2mPipe_m2sPipe_payload = counterValidAddrOneStream_s2mPipe_rData;
  assign counterValidAddrOneStream_s2mPipe_m2sPipe_ready = ((! CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready) || CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready = CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_counterOneValidStream_payload = CICC1851_validBufferOne_port2[0];
  assign CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_8 = readStage_counterOneValidStream_ready;
    if(when_Stream_l368_16) begin
      CICC1851_8 = 1'b1;
    end
  end

  assign when_Stream_l368_16 = (! readStage_counterOneValidStream_valid);
  assign readStage_counterOneValidStream_valid = CICC1851_readStage_counterOneValidStream_valid;
  assign readStage_counterOneValidStream_payload = CICC1851_readStage_counterOneValidStream_payload_2;
  assign mainValidAddrTwoStream_ready = (! mainValidAddrTwoStream_rValid);
  assign mainValidAddrTwoStream_s2mPipe_valid = (mainValidAddrTwoStream_valid || mainValidAddrTwoStream_rValid);
  assign mainValidAddrTwoStream_s2mPipe_payload = (mainValidAddrTwoStream_rValid ? mainValidAddrTwoStream_rData : mainValidAddrTwoStream_payload);
  always @(*) begin
    mainValidAddrTwoStream_s2mPipe_ready = mainValidAddrTwoStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_17) begin
      mainValidAddrTwoStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_17 = (! mainValidAddrTwoStream_s2mPipe_m2sPipe_valid);
  assign mainValidAddrTwoStream_s2mPipe_m2sPipe_valid = mainValidAddrTwoStream_s2mPipe_rValid;
  assign mainValidAddrTwoStream_s2mPipe_m2sPipe_payload = mainValidAddrTwoStream_s2mPipe_rData;
  assign mainValidAddrTwoStream_s2mPipe_m2sPipe_ready = ((! CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready) || CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready = CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_mainTwoValidStream_payload = CICC1851_validBufferTwo_port1[0];
  assign CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_9 = readStage_mainTwoValidStream_ready;
    if(when_Stream_l368_18) begin
      CICC1851_9 = 1'b1;
    end
  end

  assign when_Stream_l368_18 = (! readStage_mainTwoValidStream_valid);
  assign readStage_mainTwoValidStream_valid = CICC1851_readStage_mainTwoValidStream_valid;
  assign readStage_mainTwoValidStream_payload = CICC1851_readStage_mainTwoValidStream_payload_2;
  assign counterValidAddrTwoStream_ready = (! counterValidAddrTwoStream_rValid);
  assign counterValidAddrTwoStream_s2mPipe_valid = (counterValidAddrTwoStream_valid || counterValidAddrTwoStream_rValid);
  assign counterValidAddrTwoStream_s2mPipe_payload = (counterValidAddrTwoStream_rValid ? counterValidAddrTwoStream_rData : counterValidAddrTwoStream_payload);
  always @(*) begin
    counterValidAddrTwoStream_s2mPipe_ready = counterValidAddrTwoStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_19) begin
      counterValidAddrTwoStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_19 = (! counterValidAddrTwoStream_s2mPipe_m2sPipe_valid);
  assign counterValidAddrTwoStream_s2mPipe_m2sPipe_valid = counterValidAddrTwoStream_s2mPipe_rValid;
  assign counterValidAddrTwoStream_s2mPipe_m2sPipe_payload = counterValidAddrTwoStream_s2mPipe_rData;
  assign counterValidAddrTwoStream_s2mPipe_m2sPipe_ready = ((! CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready) || CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready = CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_counterTwoValidStream_payload = CICC1851_validBufferTwo_port2[0];
  assign CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_10 = readStage_counterTwoValidStream_ready;
    if(when_Stream_l368_20) begin
      CICC1851_10 = 1'b1;
    end
  end

  assign when_Stream_l368_20 = (! readStage_counterTwoValidStream_valid);
  assign readStage_counterTwoValidStream_valid = CICC1851_readStage_counterTwoValidStream_valid;
  assign readStage_counterTwoValidStream_payload = CICC1851_readStage_counterTwoValidStream_payload_2;
  assign mainValidAddrThreeStream_ready = (! mainValidAddrThreeStream_rValid);
  assign mainValidAddrThreeStream_s2mPipe_valid = (mainValidAddrThreeStream_valid || mainValidAddrThreeStream_rValid);
  assign mainValidAddrThreeStream_s2mPipe_payload = (mainValidAddrThreeStream_rValid ? mainValidAddrThreeStream_rData : mainValidAddrThreeStream_payload);
  always @(*) begin
    mainValidAddrThreeStream_s2mPipe_ready = mainValidAddrThreeStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_21) begin
      mainValidAddrThreeStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_21 = (! mainValidAddrThreeStream_s2mPipe_m2sPipe_valid);
  assign mainValidAddrThreeStream_s2mPipe_m2sPipe_valid = mainValidAddrThreeStream_s2mPipe_rValid;
  assign mainValidAddrThreeStream_s2mPipe_m2sPipe_payload = mainValidAddrThreeStream_s2mPipe_rData;
  assign mainValidAddrThreeStream_s2mPipe_m2sPipe_ready = ((! CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready) || CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready = CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_mainThreeValidStream_payload = CICC1851_validBufferThree_port1[0];
  assign CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_11 = readStage_mainThreeValidStream_ready;
    if(when_Stream_l368_22) begin
      CICC1851_11 = 1'b1;
    end
  end

  assign when_Stream_l368_22 = (! readStage_mainThreeValidStream_valid);
  assign readStage_mainThreeValidStream_valid = CICC1851_readStage_mainThreeValidStream_valid;
  assign readStage_mainThreeValidStream_payload = CICC1851_readStage_mainThreeValidStream_payload_2;
  assign counterValidAddrThreeStream_ready = (! counterValidAddrThreeStream_rValid);
  assign counterValidAddrThreeStream_s2mPipe_valid = (counterValidAddrThreeStream_valid || counterValidAddrThreeStream_rValid);
  assign counterValidAddrThreeStream_s2mPipe_payload = (counterValidAddrThreeStream_rValid ? counterValidAddrThreeStream_rData : counterValidAddrThreeStream_payload);
  always @(*) begin
    counterValidAddrThreeStream_s2mPipe_ready = counterValidAddrThreeStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_23) begin
      counterValidAddrThreeStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_23 = (! counterValidAddrThreeStream_s2mPipe_m2sPipe_valid);
  assign counterValidAddrThreeStream_s2mPipe_m2sPipe_valid = counterValidAddrThreeStream_s2mPipe_rValid;
  assign counterValidAddrThreeStream_s2mPipe_m2sPipe_payload = counterValidAddrThreeStream_s2mPipe_rData;
  assign counterValidAddrThreeStream_s2mPipe_m2sPipe_ready = ((! CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready) || CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready = CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_counterThreeValidStream_payload = CICC1851_validBufferThree_port2[0];
  assign CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_12 = readStage_counterThreeValidStream_ready;
    if(when_Stream_l368_24) begin
      CICC1851_12 = 1'b1;
    end
  end

  assign when_Stream_l368_24 = (! readStage_counterThreeValidStream_valid);
  assign readStage_counterThreeValidStream_valid = CICC1851_readStage_counterThreeValidStream_valid;
  assign readStage_counterThreeValidStream_payload = CICC1851_readStage_counterThreeValidStream_payload_2;
  assign controlStream_ready = (! controlStream_rValid);
  assign controlStream_s2mPipe_valid = (controlStream_valid || controlStream_rValid);
  assign controlStream_s2mPipe_payload_frameStart = (controlStream_rValid ? controlStream_rData_frameStart : controlStream_payload_frameStart);
  assign controlStream_s2mPipe_payload_rowEnd = (controlStream_rValid ? controlStream_rData_rowEnd : controlStream_payload_rowEnd);
  assign controlStream_s2mPipe_payload_pipeValid = (controlStream_rValid ? controlStream_rData_pipeValid : controlStream_payload_pipeValid);
  assign controlStream_s2mPipe_payload_firstRow = (controlStream_rValid ? controlStream_rData_firstRow : controlStream_payload_firstRow);
  assign controlStream_s2mPipe_payload_lastRow = (controlStream_rValid ? controlStream_rData_lastRow : controlStream_payload_lastRow);
  assign controlStream_s2mPipe_payload_finalResult = (controlStream_rValid ? controlStream_rData_finalResult : controlStream_payload_finalResult);
  assign controlStream_s2mPipe_payload_mainCompare = (controlStream_rValid ? controlStream_rData_mainCompare : controlStream_payload_mainCompare);
  assign controlStream_s2mPipe_payload_counterCompare = (controlStream_rValid ? controlStream_rData_counterCompare : controlStream_payload_counterCompare);
  assign controlStream_s2mPipe_payload_horizontalCompare = (controlStream_rValid ? controlStream_rData_horizontalCompare : controlStream_payload_horizontalCompare);
  assign controlStream_s2mPipe_payload_verticalCompare = (controlStream_rValid ? controlStream_rData_verticalCompare : controlStream_payload_verticalCompare);
  assign controlStream_s2mPipe_payload_mainDiff = (controlStream_rValid ? controlStream_rData_mainDiff : controlStream_payload_mainDiff);
  assign controlStream_s2mPipe_payload_counterDiff = (controlStream_rValid ? controlStream_rData_counterDiff : controlStream_payload_counterDiff);
  assign controlStream_s2mPipe_payload_horizontalDiff = (controlStream_rValid ? controlStream_rData_horizontalDiff : controlStream_payload_horizontalDiff);
  assign controlStream_s2mPipe_payload_verticalDiff = (controlStream_rValid ? controlStream_rData_verticalDiff : controlStream_payload_verticalDiff);
  assign controlStream_s2mPipe_payload_isHorizontalMin = (controlStream_rValid ? controlStream_rData_isHorizontalMin : controlStream_payload_isHorizontalMin);
  assign controlStream_s2mPipe_payload_minDiff = (controlStream_rValid ? controlStream_rData_minDiff : controlStream_payload_minDiff);
  assign controlStream_s2mPipe_payload_currentPosition = (controlStream_rValid ? controlStream_rData_currentPosition : controlStream_payload_currentPosition);
  assign controlStream_s2mPipe_payload_nextPosition = (controlStream_rValid ? controlStream_rData_nextPosition : controlStream_payload_nextPosition);
  assign controlStream_s2mPipe_payload_horizontalDirectionValid = (controlStream_rValid ? controlStream_rData_horizontalDirectionValid : controlStream_payload_horizontalDirectionValid);
  assign controlStream_s2mPipe_payload_verticalDirectionValid = (controlStream_rValid ? controlStream_rData_verticalDirectionValid : controlStream_payload_verticalDirectionValid);
  assign controlStream_s2mPipe_payload_mainDirectionValid = (controlStream_rValid ? controlStream_rData_mainDirectionValid : controlStream_payload_mainDirectionValid);
  assign controlStream_s2mPipe_payload_counterDirectionValid = (controlStream_rValid ? controlStream_rData_counterDirectionValid : controlStream_payload_counterDirectionValid);
  assign controlStream_s2mPipe_payload_inValidMinDiff = (controlStream_rValid ? controlStream_rData_inValidMinDiff : controlStream_payload_inValidMinDiff);
  always @(*) begin
    controlStream_s2mPipe_ready = controlStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_25) begin
      controlStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_25 = (! controlStream_s2mPipe_m2sPipe_valid);
  assign controlStream_s2mPipe_m2sPipe_valid = controlStream_s2mPipe_rValid;
  assign controlStream_s2mPipe_m2sPipe_payload_frameStart = controlStream_s2mPipe_rData_frameStart;
  assign controlStream_s2mPipe_m2sPipe_payload_rowEnd = controlStream_s2mPipe_rData_rowEnd;
  assign controlStream_s2mPipe_m2sPipe_payload_pipeValid = controlStream_s2mPipe_rData_pipeValid;
  assign controlStream_s2mPipe_m2sPipe_payload_firstRow = controlStream_s2mPipe_rData_firstRow;
  assign controlStream_s2mPipe_m2sPipe_payload_lastRow = controlStream_s2mPipe_rData_lastRow;
  assign controlStream_s2mPipe_m2sPipe_payload_finalResult = controlStream_s2mPipe_rData_finalResult;
  assign controlStream_s2mPipe_m2sPipe_payload_mainCompare = controlStream_s2mPipe_rData_mainCompare;
  assign controlStream_s2mPipe_m2sPipe_payload_counterCompare = controlStream_s2mPipe_rData_counterCompare;
  assign controlStream_s2mPipe_m2sPipe_payload_horizontalCompare = controlStream_s2mPipe_rData_horizontalCompare;
  assign controlStream_s2mPipe_m2sPipe_payload_verticalCompare = controlStream_s2mPipe_rData_verticalCompare;
  assign controlStream_s2mPipe_m2sPipe_payload_mainDiff = controlStream_s2mPipe_rData_mainDiff;
  assign controlStream_s2mPipe_m2sPipe_payload_counterDiff = controlStream_s2mPipe_rData_counterDiff;
  assign controlStream_s2mPipe_m2sPipe_payload_horizontalDiff = controlStream_s2mPipe_rData_horizontalDiff;
  assign controlStream_s2mPipe_m2sPipe_payload_verticalDiff = controlStream_s2mPipe_rData_verticalDiff;
  assign controlStream_s2mPipe_m2sPipe_payload_isHorizontalMin = controlStream_s2mPipe_rData_isHorizontalMin;
  assign controlStream_s2mPipe_m2sPipe_payload_minDiff = controlStream_s2mPipe_rData_minDiff;
  assign controlStream_s2mPipe_m2sPipe_payload_currentPosition = controlStream_s2mPipe_rData_currentPosition;
  assign controlStream_s2mPipe_m2sPipe_payload_nextPosition = controlStream_s2mPipe_rData_nextPosition;
  assign controlStream_s2mPipe_m2sPipe_payload_horizontalDirectionValid = controlStream_s2mPipe_rData_horizontalDirectionValid;
  assign controlStream_s2mPipe_m2sPipe_payload_verticalDirectionValid = controlStream_s2mPipe_rData_verticalDirectionValid;
  assign controlStream_s2mPipe_m2sPipe_payload_mainDirectionValid = controlStream_s2mPipe_rData_mainDirectionValid;
  assign controlStream_s2mPipe_m2sPipe_payload_counterDirectionValid = controlStream_s2mPipe_rData_counterDirectionValid;
  assign controlStream_s2mPipe_m2sPipe_payload_inValidMinDiff = controlStream_s2mPipe_rData_inValidMinDiff;
  always @(*) begin
    controlStream_s2mPipe_m2sPipe_ready = controlStream_s2mPipe_m2sPipe_m2sPipe_ready;
    if(when_Stream_l368_26) begin
      controlStream_s2mPipe_m2sPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_26 = (! controlStream_s2mPipe_m2sPipe_m2sPipe_valid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_valid = controlStream_s2mPipe_m2sPipe_rValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_frameStart = controlStream_s2mPipe_m2sPipe_rData_frameStart;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_rowEnd = controlStream_s2mPipe_m2sPipe_rData_rowEnd;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_pipeValid = controlStream_s2mPipe_m2sPipe_rData_pipeValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_firstRow = controlStream_s2mPipe_m2sPipe_rData_firstRow;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_lastRow = controlStream_s2mPipe_m2sPipe_rData_lastRow;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_finalResult = controlStream_s2mPipe_m2sPipe_rData_finalResult;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainCompare = controlStream_s2mPipe_m2sPipe_rData_mainCompare;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterCompare = controlStream_s2mPipe_m2sPipe_rData_counterCompare;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_horizontalCompare = controlStream_s2mPipe_m2sPipe_rData_horizontalCompare;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_verticalCompare = controlStream_s2mPipe_m2sPipe_rData_verticalCompare;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDiff = controlStream_s2mPipe_m2sPipe_rData_mainDiff;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDiff = controlStream_s2mPipe_m2sPipe_rData_counterDiff;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_horizontalDiff = controlStream_s2mPipe_m2sPipe_rData_horizontalDiff;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_verticalDiff = controlStream_s2mPipe_m2sPipe_rData_verticalDiff;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_isHorizontalMin = controlStream_s2mPipe_m2sPipe_rData_isHorizontalMin;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_minDiff = controlStream_s2mPipe_m2sPipe_rData_minDiff;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_currentPosition = controlStream_s2mPipe_m2sPipe_rData_currentPosition;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_nextPosition = controlStream_s2mPipe_m2sPipe_rData_nextPosition;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_horizontalDirectionValid = controlStream_s2mPipe_m2sPipe_rData_horizontalDirectionValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_verticalDirectionValid = controlStream_s2mPipe_m2sPipe_rData_verticalDirectionValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDirectionValid = controlStream_s2mPipe_m2sPipe_rData_mainDirectionValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDirectionValid = controlStream_s2mPipe_m2sPipe_rData_counterDirectionValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_inValidMinDiff = controlStream_s2mPipe_m2sPipe_rData_inValidMinDiff;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_ready = (! controlStream_s2mPipe_m2sPipe_m2sPipe_rValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_valid = (controlStream_s2mPipe_m2sPipe_m2sPipe_valid || controlStream_s2mPipe_m2sPipe_m2sPipe_rValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_frameStart = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_frameStart : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_frameStart);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_rowEnd = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_rowEnd : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_rowEnd);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_pipeValid = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_pipeValid : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_pipeValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_firstRow = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_firstRow : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_firstRow);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_lastRow = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_lastRow : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_lastRow);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_finalResult = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_finalResult : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_finalResult);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainCompare = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainCompare : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainCompare);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterCompare = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterCompare : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterCompare);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_horizontalCompare = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_horizontalCompare : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_horizontalCompare);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_verticalCompare = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_verticalCompare : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_verticalCompare);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainDiff = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainDiff : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDiff);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterDiff = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterDiff : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDiff);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_horizontalDiff = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_horizontalDiff : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_horizontalDiff);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_verticalDiff = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_verticalDiff : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_verticalDiff);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_isHorizontalMin = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_isHorizontalMin : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_isHorizontalMin);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_minDiff = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_minDiff : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_minDiff);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_currentPosition = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_currentPosition : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_currentPosition);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_nextPosition = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_nextPosition : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_nextPosition);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_horizontalDirectionValid = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_horizontalDirectionValid : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_horizontalDirectionValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_verticalDirectionValid = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_verticalDirectionValid : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_verticalDirectionValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainDirectionValid = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainDirectionValid : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDirectionValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterDirectionValid = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterDirectionValid : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDirectionValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_inValidMinDiff = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_inValidMinDiff : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_inValidMinDiff);
  always @(*) begin
    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready = readStage_controlPipe_ready;
    if(when_Stream_l368_27) begin
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_27 = (! readStage_controlPipe_valid);
  assign readStage_controlPipe_valid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rValid;
  assign readStage_controlPipe_payload_frameStart = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_frameStart;
  assign readStage_controlPipe_payload_rowEnd = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_rowEnd;
  assign readStage_controlPipe_payload_pipeValid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_pipeValid;
  assign readStage_controlPipe_payload_firstRow = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_firstRow;
  assign readStage_controlPipe_payload_lastRow = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_lastRow;
  assign readStage_controlPipe_payload_finalResult = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_finalResult;
  assign readStage_controlPipe_payload_mainCompare = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainCompare;
  assign readStage_controlPipe_payload_counterCompare = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterCompare;
  assign readStage_controlPipe_payload_horizontalCompare = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_horizontalCompare;
  assign readStage_controlPipe_payload_verticalCompare = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_verticalCompare;
  assign readStage_controlPipe_payload_mainDiff = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainDiff;
  assign readStage_controlPipe_payload_counterDiff = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterDiff;
  assign readStage_controlPipe_payload_horizontalDiff = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_horizontalDiff;
  assign readStage_controlPipe_payload_verticalDiff = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_verticalDiff;
  assign readStage_controlPipe_payload_isHorizontalMin = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_isHorizontalMin;
  assign readStage_controlPipe_payload_minDiff = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_minDiff;
  assign readStage_controlPipe_payload_currentPosition = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_currentPosition;
  assign readStage_controlPipe_payload_nextPosition = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_nextPosition;
  assign readStage_controlPipe_payload_horizontalDirectionValid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_horizontalDirectionValid;
  assign readStage_controlPipe_payload_verticalDirectionValid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_verticalDirectionValid;
  assign readStage_controlPipe_payload_mainDirectionValid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainDirectionValid;
  assign readStage_controlPipe_payload_counterDirectionValid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterDirectionValid;
  assign readStage_controlPipe_payload_inValidMinDiff = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_inValidMinDiff;
  assign readStage_mainOnePixelStream_ready = (! readStage_mainOnePixelStream_rValid);
  assign readStage_mainOnePixelStream_s2mPipe_valid = (readStage_mainOnePixelStream_valid || readStage_mainOnePixelStream_rValid);
  assign readStage_mainOnePixelStream_s2mPipe_payload = (readStage_mainOnePixelStream_rValid ? readStage_mainOnePixelStream_rData : readStage_mainOnePixelStream_payload);
  always @(*) begin
    readStage_mainOnePixelStream_s2mPipe_ready = compareStage_mainOnePixelStream_ready;
    if(when_Stream_l368_28) begin
      readStage_mainOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_28 = (! compareStage_mainOnePixelStream_valid);
  assign compareStage_mainOnePixelStream_valid = readStage_mainOnePixelStream_s2mPipe_rValid;
  assign compareStage_mainOnePixelStream_payload = readStage_mainOnePixelStream_s2mPipe_rData;
  assign readStage_counterOnePixelStream_ready = (! readStage_counterOnePixelStream_rValid);
  assign readStage_counterOnePixelStream_s2mPipe_valid = (readStage_counterOnePixelStream_valid || readStage_counterOnePixelStream_rValid);
  assign readStage_counterOnePixelStream_s2mPipe_payload = (readStage_counterOnePixelStream_rValid ? readStage_counterOnePixelStream_rData : readStage_counterOnePixelStream_payload);
  always @(*) begin
    readStage_counterOnePixelStream_s2mPipe_ready = compareStage_counterOnePixelStream_ready;
    if(when_Stream_l368_29) begin
      readStage_counterOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_29 = (! compareStage_counterOnePixelStream_valid);
  assign compareStage_counterOnePixelStream_valid = readStage_counterOnePixelStream_s2mPipe_rValid;
  assign compareStage_counterOnePixelStream_payload = readStage_counterOnePixelStream_s2mPipe_rData;
  assign readStage_mainTwoPixelStream_ready = (! readStage_mainTwoPixelStream_rValid);
  assign readStage_mainTwoPixelStream_s2mPipe_valid = (readStage_mainTwoPixelStream_valid || readStage_mainTwoPixelStream_rValid);
  assign readStage_mainTwoPixelStream_s2mPipe_payload = (readStage_mainTwoPixelStream_rValid ? readStage_mainTwoPixelStream_rData : readStage_mainTwoPixelStream_payload);
  always @(*) begin
    readStage_mainTwoPixelStream_s2mPipe_ready = compareStage_mainTwoPixelStream_ready;
    if(when_Stream_l368_30) begin
      readStage_mainTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_30 = (! compareStage_mainTwoPixelStream_valid);
  assign compareStage_mainTwoPixelStream_valid = readStage_mainTwoPixelStream_s2mPipe_rValid;
  assign compareStage_mainTwoPixelStream_payload = readStage_mainTwoPixelStream_s2mPipe_rData;
  assign readStage_counterTwoPixelStream_ready = (! readStage_counterTwoPixelStream_rValid);
  assign readStage_counterTwoPixelStream_s2mPipe_valid = (readStage_counterTwoPixelStream_valid || readStage_counterTwoPixelStream_rValid);
  assign readStage_counterTwoPixelStream_s2mPipe_payload = (readStage_counterTwoPixelStream_rValid ? readStage_counterTwoPixelStream_rData : readStage_counterTwoPixelStream_payload);
  always @(*) begin
    readStage_counterTwoPixelStream_s2mPipe_ready = compareStage_counterTwoPixelStream_ready;
    if(when_Stream_l368_31) begin
      readStage_counterTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_31 = (! compareStage_counterTwoPixelStream_valid);
  assign compareStage_counterTwoPixelStream_valid = readStage_counterTwoPixelStream_s2mPipe_rValid;
  assign compareStage_counterTwoPixelStream_payload = readStage_counterTwoPixelStream_s2mPipe_rData;
  assign readStage_mainThreePixelStream_ready = (! readStage_mainThreePixelStream_rValid);
  assign readStage_mainThreePixelStream_s2mPipe_valid = (readStage_mainThreePixelStream_valid || readStage_mainThreePixelStream_rValid);
  assign readStage_mainThreePixelStream_s2mPipe_payload = (readStage_mainThreePixelStream_rValid ? readStage_mainThreePixelStream_rData : readStage_mainThreePixelStream_payload);
  always @(*) begin
    readStage_mainThreePixelStream_s2mPipe_ready = compareStage_mainThreePixelStream_ready;
    if(when_Stream_l368_32) begin
      readStage_mainThreePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_32 = (! compareStage_mainThreePixelStream_valid);
  assign compareStage_mainThreePixelStream_valid = readStage_mainThreePixelStream_s2mPipe_rValid;
  assign compareStage_mainThreePixelStream_payload = readStage_mainThreePixelStream_s2mPipe_rData;
  assign readStage_counterThreePixelStream_ready = (! readStage_counterThreePixelStream_rValid);
  assign readStage_counterThreePixelStream_s2mPipe_valid = (readStage_counterThreePixelStream_valid || readStage_counterThreePixelStream_rValid);
  assign readStage_counterThreePixelStream_s2mPipe_payload = (readStage_counterThreePixelStream_rValid ? readStage_counterThreePixelStream_rData : readStage_counterThreePixelStream_payload);
  always @(*) begin
    readStage_counterThreePixelStream_s2mPipe_ready = compareStage_counterThreePixelStream_ready;
    if(when_Stream_l368_33) begin
      readStage_counterThreePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_33 = (! compareStage_counterThreePixelStream_valid);
  assign compareStage_counterThreePixelStream_valid = readStage_counterThreePixelStream_s2mPipe_rValid;
  assign compareStage_counterThreePixelStream_payload = readStage_counterThreePixelStream_s2mPipe_rData;
  assign readStage_mainOneValidStream_ready = (! readStage_mainOneValidStream_rValid);
  assign readStage_mainOneValidStream_s2mPipe_valid = (readStage_mainOneValidStream_valid || readStage_mainOneValidStream_rValid);
  assign readStage_mainOneValidStream_s2mPipe_payload = (readStage_mainOneValidStream_rValid ? readStage_mainOneValidStream_rData : readStage_mainOneValidStream_payload);
  always @(*) begin
    readStage_mainOneValidStream_s2mPipe_ready = compareStage_mainOneValidStream_ready;
    if(when_Stream_l368_34) begin
      readStage_mainOneValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_34 = (! compareStage_mainOneValidStream_valid);
  assign compareStage_mainOneValidStream_valid = readStage_mainOneValidStream_s2mPipe_rValid;
  assign compareStage_mainOneValidStream_payload = readStage_mainOneValidStream_s2mPipe_rData;
  assign readStage_counterOneValidStream_ready = (! readStage_counterOneValidStream_rValid);
  assign readStage_counterOneValidStream_s2mPipe_valid = (readStage_counterOneValidStream_valid || readStage_counterOneValidStream_rValid);
  assign readStage_counterOneValidStream_s2mPipe_payload = (readStage_counterOneValidStream_rValid ? readStage_counterOneValidStream_rData : readStage_counterOneValidStream_payload);
  always @(*) begin
    readStage_counterOneValidStream_s2mPipe_ready = compareStage_counterOneValidStream_ready;
    if(when_Stream_l368_35) begin
      readStage_counterOneValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_35 = (! compareStage_counterOneValidStream_valid);
  assign compareStage_counterOneValidStream_valid = readStage_counterOneValidStream_s2mPipe_rValid;
  assign compareStage_counterOneValidStream_payload = readStage_counterOneValidStream_s2mPipe_rData;
  assign readStage_mainTwoValidStream_ready = (! readStage_mainTwoValidStream_rValid);
  assign readStage_mainTwoValidStream_s2mPipe_valid = (readStage_mainTwoValidStream_valid || readStage_mainTwoValidStream_rValid);
  assign readStage_mainTwoValidStream_s2mPipe_payload = (readStage_mainTwoValidStream_rValid ? readStage_mainTwoValidStream_rData : readStage_mainTwoValidStream_payload);
  always @(*) begin
    readStage_mainTwoValidStream_s2mPipe_ready = compareStage_mainTwoValidStream_ready;
    if(when_Stream_l368_36) begin
      readStage_mainTwoValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_36 = (! compareStage_mainTwoValidStream_valid);
  assign compareStage_mainTwoValidStream_valid = readStage_mainTwoValidStream_s2mPipe_rValid;
  assign compareStage_mainTwoValidStream_payload = readStage_mainTwoValidStream_s2mPipe_rData;
  assign readStage_counterTwoValidStream_ready = (! readStage_counterTwoValidStream_rValid);
  assign readStage_counterTwoValidStream_s2mPipe_valid = (readStage_counterTwoValidStream_valid || readStage_counterTwoValidStream_rValid);
  assign readStage_counterTwoValidStream_s2mPipe_payload = (readStage_counterTwoValidStream_rValid ? readStage_counterTwoValidStream_rData : readStage_counterTwoValidStream_payload);
  always @(*) begin
    readStage_counterTwoValidStream_s2mPipe_ready = compareStage_counterTwoValidStream_ready;
    if(when_Stream_l368_37) begin
      readStage_counterTwoValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_37 = (! compareStage_counterTwoValidStream_valid);
  assign compareStage_counterTwoValidStream_valid = readStage_counterTwoValidStream_s2mPipe_rValid;
  assign compareStage_counterTwoValidStream_payload = readStage_counterTwoValidStream_s2mPipe_rData;
  assign readStage_mainThreeValidStream_ready = (! readStage_mainThreeValidStream_rValid);
  assign readStage_mainThreeValidStream_s2mPipe_valid = (readStage_mainThreeValidStream_valid || readStage_mainThreeValidStream_rValid);
  assign readStage_mainThreeValidStream_s2mPipe_payload = (readStage_mainThreeValidStream_rValid ? readStage_mainThreeValidStream_rData : readStage_mainThreeValidStream_payload);
  always @(*) begin
    readStage_mainThreeValidStream_s2mPipe_ready = compareStage_mainThreeValidStream_ready;
    if(when_Stream_l368_38) begin
      readStage_mainThreeValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_38 = (! compareStage_mainThreeValidStream_valid);
  assign compareStage_mainThreeValidStream_valid = readStage_mainThreeValidStream_s2mPipe_rValid;
  assign compareStage_mainThreeValidStream_payload = readStage_mainThreeValidStream_s2mPipe_rData;
  assign readStage_counterThreeValidStream_ready = (! readStage_counterThreeValidStream_rValid);
  assign readStage_counterThreeValidStream_s2mPipe_valid = (readStage_counterThreeValidStream_valid || readStage_counterThreeValidStream_rValid);
  assign readStage_counterThreeValidStream_s2mPipe_payload = (readStage_counterThreeValidStream_rValid ? readStage_counterThreeValidStream_rData : readStage_counterThreeValidStream_payload);
  always @(*) begin
    readStage_counterThreeValidStream_s2mPipe_ready = compareStage_counterThreeValidStream_ready;
    if(when_Stream_l368_39) begin
      readStage_counterThreeValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_39 = (! compareStage_counterThreeValidStream_valid);
  assign compareStage_counterThreeValidStream_valid = readStage_counterThreeValidStream_s2mPipe_rValid;
  assign compareStage_counterThreeValidStream_payload = readStage_counterThreeValidStream_s2mPipe_rData;
  always @(*) begin
    CICC1851_readStage_controlPipe_translated_payload_mainCompare = readStage_controlPipe_payload_mainCompare;
    if(!readStage_controlPipe_payload_finalResult) begin
      if(when_SuperResolutionPart3_l415) begin
        if(when_SuperResolutionPart3_l422) begin
          if(readStage_controlPipe_payload_firstRow) begin
            if(when_SuperResolutionPart3_l432) begin
              CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l449) begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l463) begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
              end
            end
          end
        end else begin
          if(readStage_controlPipe_payload_lastRow) begin
            if(when_SuperResolutionPart3_l477) begin
              CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
            end
          end else begin
            if(when_SuperResolutionPart3_l490) begin
              CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
            end
          end
        end
      end else begin
        if(when_SuperResolutionPart3_l496) begin
          if(when_SuperResolutionPart3_l502) begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l511) begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l524) begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
              end
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l539) begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l552) begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
              end
            end
          end
        end else begin
          if(when_SuperResolutionPart3_l564) begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l573) begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l586) begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
              end
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l601) begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l614) begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
              end
            end
          end
        end
      end
    end
  end

  always @(*) begin
    CICC1851_readStage_controlPipe_translated_payload_counterCompare = readStage_controlPipe_payload_counterCompare;
    if(!readStage_controlPipe_payload_finalResult) begin
      if(when_SuperResolutionPart3_l415) begin
        if(when_SuperResolutionPart3_l422) begin
          if(readStage_controlPipe_payload_firstRow) begin
            if(when_SuperResolutionPart3_l432) begin
              CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l449) begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l465) begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
              end
            end
          end
        end else begin
          if(readStage_controlPipe_payload_lastRow) begin
            if(when_SuperResolutionPart3_l477) begin
              CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
            end
          end else begin
            if(when_SuperResolutionPart3_l492) begin
              CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
            end
          end
        end
      end else begin
        if(when_SuperResolutionPart3_l496) begin
          if(when_SuperResolutionPart3_l502) begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l511) begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l526) begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
              end
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l539) begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l554) begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
              end
            end
          end
        end else begin
          if(when_SuperResolutionPart3_l564) begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l573) begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l588) begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
              end
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l601) begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l616) begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
              end
            end
          end
        end
      end
    end
  end

  always @(*) begin
    CICC1851_readStage_controlPipe_translated_payload_horizontalCompare = readStage_controlPipe_payload_horizontalCompare;
    if(!readStage_controlPipe_payload_finalResult) begin
      if(when_SuperResolutionPart3_l415) begin
        if(when_SuperResolutionPart3_l419) begin
          CICC1851_readStage_controlPipe_translated_payload_horizontalCompare = 1'b1;
        end else begin
          CICC1851_readStage_controlPipe_translated_payload_horizontalCompare = 1'b0;
        end
      end else begin
        if(when_SuperResolutionPart3_l496) begin
          if(when_SuperResolutionPart3_l500) begin
            CICC1851_readStage_controlPipe_translated_payload_horizontalCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_horizontalCompare = 1'b0;
          end
        end else begin
          if(when_SuperResolutionPart3_l562) begin
            CICC1851_readStage_controlPipe_translated_payload_horizontalCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_horizontalCompare = 1'b0;
          end
        end
      end
    end
  end

  always @(*) begin
    CICC1851_readStage_controlPipe_translated_payload_verticalCompare = readStage_controlPipe_payload_verticalCompare;
    if(readStage_controlPipe_payload_finalResult) begin
      if(when_SuperResolutionPart3_l342) begin
        CICC1851_readStage_controlPipe_translated_payload_verticalCompare = 1'b1;
      end else begin
        if(when_SuperResolutionPart3_l344) begin
          if(when_SuperResolutionPart3_l345) begin
            CICC1851_readStage_controlPipe_translated_payload_verticalCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_verticalCompare = 1'b0;
          end
        end else begin
          if(when_SuperResolutionPart3_l347) begin
            if(when_SuperResolutionPart3_l348) begin
              CICC1851_readStage_controlPipe_translated_payload_verticalCompare = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_verticalCompare = 1'b0;
            end
          end else begin
            if(when_SuperResolutionPart3_l351) begin
              CICC1851_readStage_controlPipe_translated_payload_verticalCompare = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_verticalCompare = 1'b0;
            end
          end
        end
      end
    end
  end

  always @(*) begin
    CICC1851_readStage_controlPipe_translated_payload_horizontalDirectionValid = readStage_controlPipe_payload_horizontalDirectionValid;
    if(!readStage_controlPipe_payload_finalResult) begin
      if(when_SuperResolutionPart3_l415) begin
        if(when_SuperResolutionPart3_l416) begin
          CICC1851_readStage_controlPipe_translated_payload_horizontalDirectionValid = 1'b1;
        end else begin
          CICC1851_readStage_controlPipe_translated_payload_horizontalDirectionValid = 1'b0;
        end
      end else begin
        if(when_SuperResolutionPart3_l496) begin
          if(when_SuperResolutionPart3_l497) begin
            CICC1851_readStage_controlPipe_translated_payload_horizontalDirectionValid = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_horizontalDirectionValid = 1'b0;
          end
        end else begin
          if(when_SuperResolutionPart3_l559) begin
            CICC1851_readStage_controlPipe_translated_payload_horizontalDirectionValid = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_horizontalDirectionValid = 1'b0;
          end
        end
      end
    end
  end

  always @(*) begin
    CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = readStage_controlPipe_payload_verticalDirectionValid;
    if(readStage_controlPipe_payload_finalResult) begin
      if(when_SuperResolutionPart3_l356) begin
        if(when_SuperResolutionPart3_l357) begin
          if(readStage_controlPipe_payload_firstRow) begin
            if(readStage_mainTwoValidStream_payload) begin
              CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b0;
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(readStage_mainThreeValidStream_payload) begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l365) begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b0;
              end
            end
          end
        end else begin
          if(readStage_controlPipe_payload_lastRow) begin
            if(readStage_mainTwoValidStream_payload) begin
              CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b0;
            end
          end else begin
            if(when_SuperResolutionPart3_l373) begin
              CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b0;
            end
          end
        end
      end else begin
        if(when_SuperResolutionPart3_l377) begin
          if(when_SuperResolutionPart3_l378) begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(readStage_mainThreeValidStream_payload) begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l383) begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b0;
              end
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(readStage_mainOneValidStream_payload) begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l391) begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b0;
              end
            end
          end
        end else begin
          if(when_SuperResolutionPart3_l396) begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(readStage_mainTwoValidStream_payload) begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l401) begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b0;
              end
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(readStage_mainOneValidStream_payload) begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l409) begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b0;
              end
            end
          end
        end
      end
    end
  end

  always @(*) begin
    CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = readStage_controlPipe_payload_mainDirectionValid;
    if(!readStage_controlPipe_payload_finalResult) begin
      if(when_SuperResolutionPart3_l415) begin
        if(when_SuperResolutionPart3_l422) begin
          if(readStage_controlPipe_payload_firstRow) begin
            if(when_SuperResolutionPart3_l424) begin
              CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b0;
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l441) begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l458) begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b0;
              end
            end
          end
        end else begin
          if(readStage_controlPipe_payload_lastRow) begin
            if(when_SuperResolutionPart3_l470) begin
              CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b0;
            end
          end else begin
            if(when_SuperResolutionPart3_l485) begin
              CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b0;
            end
          end
        end
      end else begin
        if(when_SuperResolutionPart3_l496) begin
          if(when_SuperResolutionPart3_l502) begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l504) begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l519) begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b0;
              end
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l531) begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l547) begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b0;
              end
            end
          end
        end else begin
          if(when_SuperResolutionPart3_l564) begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l566) begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l581) begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b0;
              end
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l593) begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l609) begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b0;
              end
            end
          end
        end
      end
    end
  end

  always @(*) begin
    CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = readStage_controlPipe_payload_counterDirectionValid;
    if(!readStage_controlPipe_payload_finalResult) begin
      if(when_SuperResolutionPart3_l415) begin
        if(when_SuperResolutionPart3_l422) begin
          if(readStage_controlPipe_payload_firstRow) begin
            if(when_SuperResolutionPart3_l424) begin
              CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b0;
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l441) begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l460) begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b0;
              end
            end
          end
        end else begin
          if(readStage_controlPipe_payload_lastRow) begin
            if(when_SuperResolutionPart3_l470) begin
              CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b0;
            end
          end else begin
            if(when_SuperResolutionPart3_l487) begin
              CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b0;
            end
          end
        end
      end else begin
        if(when_SuperResolutionPart3_l496) begin
          if(when_SuperResolutionPart3_l502) begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l504) begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l521) begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b0;
              end
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l531) begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l549) begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b0;
              end
            end
          end
        end else begin
          if(when_SuperResolutionPart3_l564) begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l566) begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l583) begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b0;
              end
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l593) begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l611) begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b0;
              end
            end
          end
        end
      end
    end
  end

  assign when_SuperResolutionPart3_l342 = (readStage_controlPipe_payload_firstRow || readStage_controlPipe_payload_lastRow);
  assign when_SuperResolutionPart3_l344 = (readStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l345 = (readStage_mainThreePixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart3_l348 = (readStage_mainThreePixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart3_l351 = (readStage_mainTwoPixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart3_l347 = (readStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l356 = (readStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l357 = (readStage_controlPipe_payload_nextPosition == 2'b01);
  assign when_SuperResolutionPart3_l365 = (readStage_mainTwoValidStream_payload && readStage_mainThreeValidStream_payload);
  assign when_SuperResolutionPart3_l373 = (readStage_mainTwoValidStream_payload && readStage_mainThreeValidStream_payload);
  assign when_SuperResolutionPart3_l378 = (readStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l383 = (readStage_mainOneValidStream_payload && readStage_mainThreeValidStream_payload);
  assign when_SuperResolutionPart3_l391 = (readStage_mainOneValidStream_payload && readStage_mainThreeValidStream_payload);
  assign when_SuperResolutionPart3_l396 = (readStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l401 = (readStage_mainOneValidStream_payload && readStage_mainTwoValidStream_payload);
  assign when_SuperResolutionPart3_l409 = (readStage_mainOneValidStream_payload && readStage_mainTwoValidStream_payload);
  assign when_SuperResolutionPart3_l377 = (readStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l415 = (readStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l416 = (readStage_mainOneValidStream_payload && readStage_counterOneValidStream_payload);
  assign when_SuperResolutionPart3_l419 = (readStage_counterOnePixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart3_l422 = (readStage_controlPipe_payload_nextPosition == 2'b01);
  assign when_SuperResolutionPart3_l424 = (readStage_mainTwoValidStream_payload && readStage_counterTwoValidStream_payload);
  assign when_SuperResolutionPart3_l432 = (readStage_counterTwoPixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart3_l441 = (readStage_mainThreeValidStream_payload && readStage_counterThreeValidStream_payload);
  assign when_SuperResolutionPart3_l449 = (readStage_counterThreePixelStream_payload <= readStage_mainThreePixelStream_payload);
  assign when_SuperResolutionPart3_l458 = (readStage_mainThreeValidStream_payload && readStage_counterTwoValidStream_payload);
  assign when_SuperResolutionPart3_l460 = (readStage_mainTwoValidStream_payload && readStage_counterThreeValidStream_payload);
  assign when_SuperResolutionPart3_l463 = (readStage_counterTwoPixelStream_payload <= readStage_mainThreePixelStream_payload);
  assign when_SuperResolutionPart3_l465 = (readStage_counterThreePixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart3_l470 = (readStage_mainTwoValidStream_payload && readStage_counterTwoValidStream_payload);
  assign when_SuperResolutionPart3_l477 = (readStage_counterTwoPixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart3_l485 = (readStage_mainTwoValidStream_payload && readStage_counterThreeValidStream_payload);
  assign when_SuperResolutionPart3_l487 = (readStage_mainThreeValidStream_payload && readStage_counterTwoValidStream_payload);
  assign when_SuperResolutionPart3_l490 = (readStage_counterThreePixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart3_l492 = (readStage_counterTwoPixelStream_payload <= readStage_mainThreePixelStream_payload);
  assign when_SuperResolutionPart3_l497 = (readStage_mainTwoValidStream_payload && readStage_counterTwoValidStream_payload);
  assign when_SuperResolutionPart3_l500 = (readStage_counterTwoPixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart3_l502 = (readStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l504 = (readStage_mainThreeValidStream_payload && readStage_counterThreeValidStream_payload);
  assign when_SuperResolutionPart3_l511 = (readStage_counterThreePixelStream_payload <= readStage_mainThreePixelStream_payload);
  assign when_SuperResolutionPart3_l519 = (readStage_mainThreeValidStream_payload && readStage_counterOneValidStream_payload);
  assign when_SuperResolutionPart3_l521 = (readStage_mainOneValidStream_payload && readStage_counterThreeValidStream_payload);
  assign when_SuperResolutionPart3_l524 = (readStage_counterOnePixelStream_payload <= readStage_mainThreePixelStream_payload);
  assign when_SuperResolutionPart3_l526 = (readStage_counterThreePixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart3_l531 = (readStage_mainOneValidStream_payload && readStage_counterOneValidStream_payload);
  assign when_SuperResolutionPart3_l539 = (readStage_counterOnePixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart3_l547 = (readStage_mainOneValidStream_payload && readStage_counterThreeValidStream_payload);
  assign when_SuperResolutionPart3_l549 = (readStage_mainThreeValidStream_payload && readStage_counterOneValidStream_payload);
  assign when_SuperResolutionPart3_l552 = (readStage_counterThreePixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart3_l554 = (readStage_counterOnePixelStream_payload <= readStage_mainThreePixelStream_payload);
  assign when_SuperResolutionPart3_l559 = (readStage_mainThreeValidStream_payload && readStage_counterThreeValidStream_payload);
  assign when_SuperResolutionPart3_l562 = (readStage_counterThreePixelStream_payload <= readStage_mainThreePixelStream_payload);
  assign when_SuperResolutionPart3_l564 = (readStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l566 = (readStage_mainTwoValidStream_payload && readStage_counterTwoValidStream_payload);
  assign when_SuperResolutionPart3_l573 = (readStage_counterTwoPixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart3_l581 = (readStage_mainTwoValidStream_payload && readStage_counterOneValidStream_payload);
  assign when_SuperResolutionPart3_l583 = (readStage_mainOneValidStream_payload && readStage_counterTwoValidStream_payload);
  assign when_SuperResolutionPart3_l586 = (readStage_counterOnePixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart3_l588 = (readStage_counterTwoPixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart3_l593 = (readStage_mainOneValidStream_payload && readStage_counterOneValidStream_payload);
  assign when_SuperResolutionPart3_l601 = (readStage_counterOnePixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart3_l609 = (readStage_mainOneValidStream_payload && readStage_counterTwoValidStream_payload);
  assign when_SuperResolutionPart3_l611 = (readStage_mainTwoValidStream_payload && readStage_counterOneValidStream_payload);
  assign when_SuperResolutionPart3_l614 = (readStage_counterTwoPixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart3_l616 = (readStage_counterOnePixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart3_l496 = (readStage_controlPipe_payload_currentPosition == 2'b01);
  assign readStage_controlPipe_translated_valid = readStage_controlPipe_valid;
  assign readStage_controlPipe_ready = readStage_controlPipe_translated_ready;
  assign readStage_controlPipe_translated_payload_frameStart = readStage_controlPipe_payload_frameStart;
  assign readStage_controlPipe_translated_payload_rowEnd = readStage_controlPipe_payload_rowEnd;
  assign readStage_controlPipe_translated_payload_pipeValid = readStage_controlPipe_payload_pipeValid;
  assign readStage_controlPipe_translated_payload_firstRow = readStage_controlPipe_payload_firstRow;
  assign readStage_controlPipe_translated_payload_lastRow = readStage_controlPipe_payload_lastRow;
  assign readStage_controlPipe_translated_payload_finalResult = readStage_controlPipe_payload_finalResult;
  assign readStage_controlPipe_translated_payload_mainCompare = CICC1851_readStage_controlPipe_translated_payload_mainCompare;
  assign readStage_controlPipe_translated_payload_counterCompare = CICC1851_readStage_controlPipe_translated_payload_counterCompare;
  assign readStage_controlPipe_translated_payload_horizontalCompare = CICC1851_readStage_controlPipe_translated_payload_horizontalCompare;
  assign readStage_controlPipe_translated_payload_verticalCompare = CICC1851_readStage_controlPipe_translated_payload_verticalCompare;
  assign readStage_controlPipe_translated_payload_mainDiff = readStage_controlPipe_payload_mainDiff;
  assign readStage_controlPipe_translated_payload_counterDiff = readStage_controlPipe_payload_counterDiff;
  assign readStage_controlPipe_translated_payload_horizontalDiff = readStage_controlPipe_payload_horizontalDiff;
  assign readStage_controlPipe_translated_payload_verticalDiff = readStage_controlPipe_payload_verticalDiff;
  assign readStage_controlPipe_translated_payload_isHorizontalMin = readStage_controlPipe_payload_isHorizontalMin;
  assign readStage_controlPipe_translated_payload_minDiff = readStage_controlPipe_payload_minDiff;
  assign readStage_controlPipe_translated_payload_currentPosition = readStage_controlPipe_payload_currentPosition;
  assign readStage_controlPipe_translated_payload_nextPosition = readStage_controlPipe_payload_nextPosition;
  assign readStage_controlPipe_translated_payload_horizontalDirectionValid = CICC1851_readStage_controlPipe_translated_payload_horizontalDirectionValid;
  assign readStage_controlPipe_translated_payload_verticalDirectionValid = CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid;
  assign readStage_controlPipe_translated_payload_mainDirectionValid = CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid;
  assign readStage_controlPipe_translated_payload_counterDirectionValid = CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid;
  assign readStage_controlPipe_translated_payload_inValidMinDiff = readStage_controlPipe_payload_inValidMinDiff;
  assign readStage_controlPipe_translated_ready = (! readStage_controlPipe_translated_rValid);
  assign readStage_controlPipe_translated_s2mPipe_valid = (readStage_controlPipe_translated_valid || readStage_controlPipe_translated_rValid);
  assign readStage_controlPipe_translated_s2mPipe_payload_frameStart = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_frameStart : readStage_controlPipe_translated_payload_frameStart);
  assign readStage_controlPipe_translated_s2mPipe_payload_rowEnd = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_rowEnd : readStage_controlPipe_translated_payload_rowEnd);
  assign readStage_controlPipe_translated_s2mPipe_payload_pipeValid = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_pipeValid : readStage_controlPipe_translated_payload_pipeValid);
  assign readStage_controlPipe_translated_s2mPipe_payload_firstRow = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_firstRow : readStage_controlPipe_translated_payload_firstRow);
  assign readStage_controlPipe_translated_s2mPipe_payload_lastRow = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_lastRow : readStage_controlPipe_translated_payload_lastRow);
  assign readStage_controlPipe_translated_s2mPipe_payload_finalResult = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_finalResult : readStage_controlPipe_translated_payload_finalResult);
  assign readStage_controlPipe_translated_s2mPipe_payload_mainCompare = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_mainCompare : readStage_controlPipe_translated_payload_mainCompare);
  assign readStage_controlPipe_translated_s2mPipe_payload_counterCompare = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_counterCompare : readStage_controlPipe_translated_payload_counterCompare);
  assign readStage_controlPipe_translated_s2mPipe_payload_horizontalCompare = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_horizontalCompare : readStage_controlPipe_translated_payload_horizontalCompare);
  assign readStage_controlPipe_translated_s2mPipe_payload_verticalCompare = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_verticalCompare : readStage_controlPipe_translated_payload_verticalCompare);
  assign readStage_controlPipe_translated_s2mPipe_payload_mainDiff = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_mainDiff : readStage_controlPipe_translated_payload_mainDiff);
  assign readStage_controlPipe_translated_s2mPipe_payload_counterDiff = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_counterDiff : readStage_controlPipe_translated_payload_counterDiff);
  assign readStage_controlPipe_translated_s2mPipe_payload_horizontalDiff = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_horizontalDiff : readStage_controlPipe_translated_payload_horizontalDiff);
  assign readStage_controlPipe_translated_s2mPipe_payload_verticalDiff = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_verticalDiff : readStage_controlPipe_translated_payload_verticalDiff);
  assign readStage_controlPipe_translated_s2mPipe_payload_isHorizontalMin = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_isHorizontalMin : readStage_controlPipe_translated_payload_isHorizontalMin);
  assign readStage_controlPipe_translated_s2mPipe_payload_minDiff = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_minDiff : readStage_controlPipe_translated_payload_minDiff);
  assign readStage_controlPipe_translated_s2mPipe_payload_currentPosition = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_currentPosition : readStage_controlPipe_translated_payload_currentPosition);
  assign readStage_controlPipe_translated_s2mPipe_payload_nextPosition = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_nextPosition : readStage_controlPipe_translated_payload_nextPosition);
  assign readStage_controlPipe_translated_s2mPipe_payload_horizontalDirectionValid = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_horizontalDirectionValid : readStage_controlPipe_translated_payload_horizontalDirectionValid);
  assign readStage_controlPipe_translated_s2mPipe_payload_verticalDirectionValid = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_verticalDirectionValid : readStage_controlPipe_translated_payload_verticalDirectionValid);
  assign readStage_controlPipe_translated_s2mPipe_payload_mainDirectionValid = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_mainDirectionValid : readStage_controlPipe_translated_payload_mainDirectionValid);
  assign readStage_controlPipe_translated_s2mPipe_payload_counterDirectionValid = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_counterDirectionValid : readStage_controlPipe_translated_payload_counterDirectionValid);
  assign readStage_controlPipe_translated_s2mPipe_payload_inValidMinDiff = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_inValidMinDiff : readStage_controlPipe_translated_payload_inValidMinDiff);
  always @(*) begin
    readStage_controlPipe_translated_s2mPipe_ready = compareStage_controlPipe_ready;
    if(when_Stream_l368_40) begin
      readStage_controlPipe_translated_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_40 = (! compareStage_controlPipe_valid);
  assign compareStage_controlPipe_valid = readStage_controlPipe_translated_s2mPipe_rValid;
  assign compareStage_controlPipe_payload_frameStart = readStage_controlPipe_translated_s2mPipe_rData_frameStart;
  assign compareStage_controlPipe_payload_rowEnd = readStage_controlPipe_translated_s2mPipe_rData_rowEnd;
  assign compareStage_controlPipe_payload_pipeValid = readStage_controlPipe_translated_s2mPipe_rData_pipeValid;
  assign compareStage_controlPipe_payload_firstRow = readStage_controlPipe_translated_s2mPipe_rData_firstRow;
  assign compareStage_controlPipe_payload_lastRow = readStage_controlPipe_translated_s2mPipe_rData_lastRow;
  assign compareStage_controlPipe_payload_finalResult = readStage_controlPipe_translated_s2mPipe_rData_finalResult;
  assign compareStage_controlPipe_payload_mainCompare = readStage_controlPipe_translated_s2mPipe_rData_mainCompare;
  assign compareStage_controlPipe_payload_counterCompare = readStage_controlPipe_translated_s2mPipe_rData_counterCompare;
  assign compareStage_controlPipe_payload_horizontalCompare = readStage_controlPipe_translated_s2mPipe_rData_horizontalCompare;
  assign compareStage_controlPipe_payload_verticalCompare = readStage_controlPipe_translated_s2mPipe_rData_verticalCompare;
  assign compareStage_controlPipe_payload_mainDiff = readStage_controlPipe_translated_s2mPipe_rData_mainDiff;
  assign compareStage_controlPipe_payload_counterDiff = readStage_controlPipe_translated_s2mPipe_rData_counterDiff;
  assign compareStage_controlPipe_payload_horizontalDiff = readStage_controlPipe_translated_s2mPipe_rData_horizontalDiff;
  assign compareStage_controlPipe_payload_verticalDiff = readStage_controlPipe_translated_s2mPipe_rData_verticalDiff;
  assign compareStage_controlPipe_payload_isHorizontalMin = readStage_controlPipe_translated_s2mPipe_rData_isHorizontalMin;
  assign compareStage_controlPipe_payload_minDiff = readStage_controlPipe_translated_s2mPipe_rData_minDiff;
  assign compareStage_controlPipe_payload_currentPosition = readStage_controlPipe_translated_s2mPipe_rData_currentPosition;
  assign compareStage_controlPipe_payload_nextPosition = readStage_controlPipe_translated_s2mPipe_rData_nextPosition;
  assign compareStage_controlPipe_payload_horizontalDirectionValid = readStage_controlPipe_translated_s2mPipe_rData_horizontalDirectionValid;
  assign compareStage_controlPipe_payload_verticalDirectionValid = readStage_controlPipe_translated_s2mPipe_rData_verticalDirectionValid;
  assign compareStage_controlPipe_payload_mainDirectionValid = readStage_controlPipe_translated_s2mPipe_rData_mainDirectionValid;
  assign compareStage_controlPipe_payload_counterDirectionValid = readStage_controlPipe_translated_s2mPipe_rData_counterDirectionValid;
  assign compareStage_controlPipe_payload_inValidMinDiff = readStage_controlPipe_translated_s2mPipe_rData_inValidMinDiff;
  assign compareStage_mainOnePixelStream_ready = (! compareStage_mainOnePixelStream_rValid);
  assign compareStage_mainOnePixelStream_s2mPipe_valid = (compareStage_mainOnePixelStream_valid || compareStage_mainOnePixelStream_rValid);
  assign compareStage_mainOnePixelStream_s2mPipe_payload = (compareStage_mainOnePixelStream_rValid ? compareStage_mainOnePixelStream_rData : compareStage_mainOnePixelStream_payload);
  always @(*) begin
    compareStage_mainOnePixelStream_s2mPipe_ready = diffStage_mainOnePixelStream_ready;
    if(when_Stream_l368_41) begin
      compareStage_mainOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_41 = (! diffStage_mainOnePixelStream_valid);
  assign diffStage_mainOnePixelStream_valid = compareStage_mainOnePixelStream_s2mPipe_rValid;
  assign diffStage_mainOnePixelStream_payload = compareStage_mainOnePixelStream_s2mPipe_rData;
  assign compareStage_counterOnePixelStream_ready = (! compareStage_counterOnePixelStream_rValid);
  assign compareStage_counterOnePixelStream_s2mPipe_valid = (compareStage_counterOnePixelStream_valid || compareStage_counterOnePixelStream_rValid);
  assign compareStage_counterOnePixelStream_s2mPipe_payload = (compareStage_counterOnePixelStream_rValid ? compareStage_counterOnePixelStream_rData : compareStage_counterOnePixelStream_payload);
  always @(*) begin
    compareStage_counterOnePixelStream_s2mPipe_ready = diffStage_counterOnePixelStream_ready;
    if(when_Stream_l368_42) begin
      compareStage_counterOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_42 = (! diffStage_counterOnePixelStream_valid);
  assign diffStage_counterOnePixelStream_valid = compareStage_counterOnePixelStream_s2mPipe_rValid;
  assign diffStage_counterOnePixelStream_payload = compareStage_counterOnePixelStream_s2mPipe_rData;
  assign compareStage_mainTwoPixelStream_ready = (! compareStage_mainTwoPixelStream_rValid);
  assign compareStage_mainTwoPixelStream_s2mPipe_valid = (compareStage_mainTwoPixelStream_valid || compareStage_mainTwoPixelStream_rValid);
  assign compareStage_mainTwoPixelStream_s2mPipe_payload = (compareStage_mainTwoPixelStream_rValid ? compareStage_mainTwoPixelStream_rData : compareStage_mainTwoPixelStream_payload);
  always @(*) begin
    compareStage_mainTwoPixelStream_s2mPipe_ready = diffStage_mainTwoPixelStream_ready;
    if(when_Stream_l368_43) begin
      compareStage_mainTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_43 = (! diffStage_mainTwoPixelStream_valid);
  assign diffStage_mainTwoPixelStream_valid = compareStage_mainTwoPixelStream_s2mPipe_rValid;
  assign diffStage_mainTwoPixelStream_payload = compareStage_mainTwoPixelStream_s2mPipe_rData;
  assign compareStage_counterTwoPixelStream_ready = (! compareStage_counterTwoPixelStream_rValid);
  assign compareStage_counterTwoPixelStream_s2mPipe_valid = (compareStage_counterTwoPixelStream_valid || compareStage_counterTwoPixelStream_rValid);
  assign compareStage_counterTwoPixelStream_s2mPipe_payload = (compareStage_counterTwoPixelStream_rValid ? compareStage_counterTwoPixelStream_rData : compareStage_counterTwoPixelStream_payload);
  always @(*) begin
    compareStage_counterTwoPixelStream_s2mPipe_ready = diffStage_counterTwoPixelStream_ready;
    if(when_Stream_l368_44) begin
      compareStage_counterTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_44 = (! diffStage_counterTwoPixelStream_valid);
  assign diffStage_counterTwoPixelStream_valid = compareStage_counterTwoPixelStream_s2mPipe_rValid;
  assign diffStage_counterTwoPixelStream_payload = compareStage_counterTwoPixelStream_s2mPipe_rData;
  assign compareStage_mainThreePixelStream_ready = (! compareStage_mainThreePixelStream_rValid);
  assign compareStage_mainThreePixelStream_s2mPipe_valid = (compareStage_mainThreePixelStream_valid || compareStage_mainThreePixelStream_rValid);
  assign compareStage_mainThreePixelStream_s2mPipe_payload = (compareStage_mainThreePixelStream_rValid ? compareStage_mainThreePixelStream_rData : compareStage_mainThreePixelStream_payload);
  always @(*) begin
    compareStage_mainThreePixelStream_s2mPipe_ready = diffStage_mainThreePixelStream_ready;
    if(when_Stream_l368_45) begin
      compareStage_mainThreePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_45 = (! diffStage_mainThreePixelStream_valid);
  assign diffStage_mainThreePixelStream_valid = compareStage_mainThreePixelStream_s2mPipe_rValid;
  assign diffStage_mainThreePixelStream_payload = compareStage_mainThreePixelStream_s2mPipe_rData;
  assign compareStage_counterThreePixelStream_ready = (! compareStage_counterThreePixelStream_rValid);
  assign compareStage_counterThreePixelStream_s2mPipe_valid = (compareStage_counterThreePixelStream_valid || compareStage_counterThreePixelStream_rValid);
  assign compareStage_counterThreePixelStream_s2mPipe_payload = (compareStage_counterThreePixelStream_rValid ? compareStage_counterThreePixelStream_rData : compareStage_counterThreePixelStream_payload);
  always @(*) begin
    compareStage_counterThreePixelStream_s2mPipe_ready = diffStage_counterThreePixelStream_ready;
    if(when_Stream_l368_46) begin
      compareStage_counterThreePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_46 = (! diffStage_counterThreePixelStream_valid);
  assign diffStage_counterThreePixelStream_valid = compareStage_counterThreePixelStream_s2mPipe_rValid;
  assign diffStage_counterThreePixelStream_payload = compareStage_counterThreePixelStream_s2mPipe_rData;
  assign compareStage_mainOneValidStream_ready = (! compareStage_mainOneValidStream_rValid);
  assign compareStage_mainOneValidStream_s2mPipe_valid = (compareStage_mainOneValidStream_valid || compareStage_mainOneValidStream_rValid);
  assign compareStage_mainOneValidStream_s2mPipe_payload = (compareStage_mainOneValidStream_rValid ? compareStage_mainOneValidStream_rData : compareStage_mainOneValidStream_payload);
  always @(*) begin
    compareStage_mainOneValidStream_s2mPipe_ready = diffStage_mainOneValidStream_ready;
    if(when_Stream_l368_47) begin
      compareStage_mainOneValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_47 = (! diffStage_mainOneValidStream_valid);
  assign diffStage_mainOneValidStream_valid = compareStage_mainOneValidStream_s2mPipe_rValid;
  assign diffStage_mainOneValidStream_payload = compareStage_mainOneValidStream_s2mPipe_rData;
  assign compareStage_counterOneValidStream_ready = (! compareStage_counterOneValidStream_rValid);
  assign compareStage_counterOneValidStream_s2mPipe_valid = (compareStage_counterOneValidStream_valid || compareStage_counterOneValidStream_rValid);
  assign compareStage_counterOneValidStream_s2mPipe_payload = (compareStage_counterOneValidStream_rValid ? compareStage_counterOneValidStream_rData : compareStage_counterOneValidStream_payload);
  always @(*) begin
    compareStage_counterOneValidStream_s2mPipe_ready = diffStage_counterOneValidStream_ready;
    if(when_Stream_l368_48) begin
      compareStage_counterOneValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_48 = (! diffStage_counterOneValidStream_valid);
  assign diffStage_counterOneValidStream_valid = compareStage_counterOneValidStream_s2mPipe_rValid;
  assign diffStage_counterOneValidStream_payload = compareStage_counterOneValidStream_s2mPipe_rData;
  assign compareStage_mainTwoValidStream_ready = (! compareStage_mainTwoValidStream_rValid);
  assign compareStage_mainTwoValidStream_s2mPipe_valid = (compareStage_mainTwoValidStream_valid || compareStage_mainTwoValidStream_rValid);
  assign compareStage_mainTwoValidStream_s2mPipe_payload = (compareStage_mainTwoValidStream_rValid ? compareStage_mainTwoValidStream_rData : compareStage_mainTwoValidStream_payload);
  always @(*) begin
    compareStage_mainTwoValidStream_s2mPipe_ready = diffStage_mainTwoValidStream_ready;
    if(when_Stream_l368_49) begin
      compareStage_mainTwoValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_49 = (! diffStage_mainTwoValidStream_valid);
  assign diffStage_mainTwoValidStream_valid = compareStage_mainTwoValidStream_s2mPipe_rValid;
  assign diffStage_mainTwoValidStream_payload = compareStage_mainTwoValidStream_s2mPipe_rData;
  assign compareStage_counterTwoValidStream_ready = (! compareStage_counterTwoValidStream_rValid);
  assign compareStage_counterTwoValidStream_s2mPipe_valid = (compareStage_counterTwoValidStream_valid || compareStage_counterTwoValidStream_rValid);
  assign compareStage_counterTwoValidStream_s2mPipe_payload = (compareStage_counterTwoValidStream_rValid ? compareStage_counterTwoValidStream_rData : compareStage_counterTwoValidStream_payload);
  always @(*) begin
    compareStage_counterTwoValidStream_s2mPipe_ready = diffStage_counterTwoValidStream_ready;
    if(when_Stream_l368_50) begin
      compareStage_counterTwoValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_50 = (! diffStage_counterTwoValidStream_valid);
  assign diffStage_counterTwoValidStream_valid = compareStage_counterTwoValidStream_s2mPipe_rValid;
  assign diffStage_counterTwoValidStream_payload = compareStage_counterTwoValidStream_s2mPipe_rData;
  assign compareStage_mainThreeValidStream_ready = (! compareStage_mainThreeValidStream_rValid);
  assign compareStage_mainThreeValidStream_s2mPipe_valid = (compareStage_mainThreeValidStream_valid || compareStage_mainThreeValidStream_rValid);
  assign compareStage_mainThreeValidStream_s2mPipe_payload = (compareStage_mainThreeValidStream_rValid ? compareStage_mainThreeValidStream_rData : compareStage_mainThreeValidStream_payload);
  always @(*) begin
    compareStage_mainThreeValidStream_s2mPipe_ready = diffStage_mainThreeValidStream_ready;
    if(when_Stream_l368_51) begin
      compareStage_mainThreeValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_51 = (! diffStage_mainThreeValidStream_valid);
  assign diffStage_mainThreeValidStream_valid = compareStage_mainThreeValidStream_s2mPipe_rValid;
  assign diffStage_mainThreeValidStream_payload = compareStage_mainThreeValidStream_s2mPipe_rData;
  assign compareStage_counterThreeValidStream_ready = (! compareStage_counterThreeValidStream_rValid);
  assign compareStage_counterThreeValidStream_s2mPipe_valid = (compareStage_counterThreeValidStream_valid || compareStage_counterThreeValidStream_rValid);
  assign compareStage_counterThreeValidStream_s2mPipe_payload = (compareStage_counterThreeValidStream_rValid ? compareStage_counterThreeValidStream_rData : compareStage_counterThreeValidStream_payload);
  always @(*) begin
    compareStage_counterThreeValidStream_s2mPipe_ready = diffStage_counterThreeValidStream_ready;
    if(when_Stream_l368_52) begin
      compareStage_counterThreeValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_52 = (! diffStage_counterThreeValidStream_valid);
  assign diffStage_counterThreeValidStream_valid = compareStage_counterThreeValidStream_s2mPipe_rValid;
  assign diffStage_counterThreeValidStream_payload = compareStage_counterThreeValidStream_s2mPipe_rData;
  always @(*) begin
    CICC1851_compareStage_controlPipe_translated_payload_mainDiff = compareStage_controlPipe_payload_mainDiff;
    if(!compareStage_controlPipe_payload_finalResult) begin
      if(when_SuperResolutionPart3_l661) begin
        if(when_SuperResolutionPart3_l664) begin
          if(compareStage_controlPipe_payload_firstRow) begin
            if(compareStage_controlPipe_payload_mainCompare) begin
              CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterTwoPixelStream_payload);
            end else begin
              CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainTwoPixelStream_payload);
            end
          end else begin
            if(compareStage_controlPipe_payload_lastRow) begin
              if(compareStage_controlPipe_payload_mainCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainThreePixelStream_payload - compareStage_counterThreePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterThreePixelStream_payload - compareStage_mainThreePixelStream_payload);
              end
            end else begin
              if(compareStage_controlPipe_payload_mainCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainThreePixelStream_payload - compareStage_counterTwoPixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainThreePixelStream_payload);
              end
            end
          end
        end else begin
          if(compareStage_controlPipe_payload_lastRow) begin
            if(compareStage_controlPipe_payload_mainCompare) begin
              CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterTwoPixelStream_payload);
            end else begin
              CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainTwoPixelStream_payload);
            end
          end else begin
            if(compareStage_controlPipe_payload_mainCompare) begin
              CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterThreePixelStream_payload);
            end else begin
              CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterThreePixelStream_payload - compareStage_mainTwoPixelStream_payload);
            end
          end
        end
      end else begin
        if(when_SuperResolutionPart3_l694) begin
          if(when_SuperResolutionPart3_l697) begin
            if(compareStage_controlPipe_payload_lastRow) begin
              if(compareStage_controlPipe_payload_mainCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainThreePixelStream_payload - compareStage_counterThreePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterThreePixelStream_payload - compareStage_mainThreePixelStream_payload);
              end
            end else begin
              if(compareStage_controlPipe_payload_mainCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainThreePixelStream_payload - compareStage_counterOnePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterOnePixelStream_payload - compareStage_mainThreePixelStream_payload);
              end
            end
          end else begin
            if(compareStage_controlPipe_payload_lastRow) begin
              if(compareStage_controlPipe_payload_mainCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_counterOnePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterOnePixelStream_payload - compareStage_mainOnePixelStream_payload);
              end
            end else begin
              if(compareStage_controlPipe_payload_mainCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_counterThreePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterThreePixelStream_payload - compareStage_mainOnePixelStream_payload);
              end
            end
          end
        end else begin
          if(when_SuperResolutionPart3_l725) begin
            if(compareStage_controlPipe_payload_lastRow) begin
              if(compareStage_controlPipe_payload_mainCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterTwoPixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainTwoPixelStream_payload);
              end
            end else begin
              if(compareStage_controlPipe_payload_mainCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterOnePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterOnePixelStream_payload - compareStage_mainTwoPixelStream_payload);
              end
            end
          end else begin
            if(compareStage_controlPipe_payload_lastRow) begin
              if(compareStage_controlPipe_payload_mainCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_counterOnePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterOnePixelStream_payload - compareStage_mainOnePixelStream_payload);
              end
            end else begin
              if(compareStage_controlPipe_payload_mainCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_counterTwoPixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainOnePixelStream_payload);
              end
            end
          end
        end
      end
    end
  end

  always @(*) begin
    CICC1851_compareStage_controlPipe_translated_payload_counterDiff = compareStage_controlPipe_payload_counterDiff;
    if(!compareStage_controlPipe_payload_finalResult) begin
      if(when_SuperResolutionPart3_l661) begin
        if(when_SuperResolutionPart3_l664) begin
          if(compareStage_controlPipe_payload_firstRow) begin
            if(compareStage_controlPipe_payload_counterCompare) begin
              CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterTwoPixelStream_payload);
            end else begin
              CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainTwoPixelStream_payload);
            end
          end else begin
            if(compareStage_controlPipe_payload_lastRow) begin
              if(compareStage_controlPipe_payload_counterCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_mainThreePixelStream_payload - compareStage_counterThreePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterThreePixelStream_payload - compareStage_mainThreePixelStream_payload);
              end
            end else begin
              if(compareStage_controlPipe_payload_counterCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterThreePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterThreePixelStream_payload - compareStage_mainTwoPixelStream_payload);
              end
            end
          end
        end else begin
          if(compareStage_controlPipe_payload_lastRow) begin
            if(compareStage_controlPipe_payload_counterCompare) begin
              CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterTwoPixelStream_payload);
            end else begin
              CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainTwoPixelStream_payload);
            end
          end else begin
            if(compareStage_controlPipe_payload_counterCompare) begin
              CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_mainThreePixelStream_payload - compareStage_counterTwoPixelStream_payload);
            end else begin
              CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainThreePixelStream_payload);
            end
          end
        end
      end else begin
        if(when_SuperResolutionPart3_l694) begin
          if(when_SuperResolutionPart3_l697) begin
            if(compareStage_controlPipe_payload_lastRow) begin
              if(compareStage_controlPipe_payload_counterCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_mainThreePixelStream_payload - compareStage_counterThreePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterThreePixelStream_payload - compareStage_mainThreePixelStream_payload);
              end
            end else begin
              if(compareStage_controlPipe_payload_counterCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_mainOnePixelStream_payload - compareStage_counterThreePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterThreePixelStream_payload - compareStage_mainOnePixelStream_payload);
              end
            end
          end else begin
            if(compareStage_controlPipe_payload_lastRow) begin
              if(compareStage_controlPipe_payload_counterCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_mainOnePixelStream_payload - compareStage_counterOnePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterOnePixelStream_payload - compareStage_mainOnePixelStream_payload);
              end
            end else begin
              if(compareStage_controlPipe_payload_counterCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_mainThreePixelStream_payload - compareStage_counterOnePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterOnePixelStream_payload - compareStage_mainThreePixelStream_payload);
              end
            end
          end
        end else begin
          if(when_SuperResolutionPart3_l725) begin
            if(compareStage_controlPipe_payload_lastRow) begin
              if(compareStage_controlPipe_payload_counterCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterTwoPixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainTwoPixelStream_payload);
              end
            end else begin
              if(compareStage_controlPipe_payload_counterCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_mainOnePixelStream_payload - compareStage_counterTwoPixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainOnePixelStream_payload);
              end
            end
          end else begin
            if(compareStage_controlPipe_payload_lastRow) begin
              if(compareStage_controlPipe_payload_counterCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_mainOnePixelStream_payload - compareStage_counterOnePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterOnePixelStream_payload - compareStage_mainOnePixelStream_payload);
              end
            end else begin
              if(compareStage_controlPipe_payload_counterCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterOnePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterOnePixelStream_payload - compareStage_mainTwoPixelStream_payload);
              end
            end
          end
        end
      end
    end
  end

  always @(*) begin
    CICC1851_compareStage_controlPipe_translated_payload_horizontalDiff = compareStage_controlPipe_payload_horizontalDiff;
    if(!compareStage_controlPipe_payload_finalResult) begin
      if(when_SuperResolutionPart3_l661) begin
        if(compareStage_controlPipe_payload_horizontalCompare) begin
          CICC1851_compareStage_controlPipe_translated_payload_horizontalDiff = (compareStage_mainOnePixelStream_payload - compareStage_counterOnePixelStream_payload);
        end else begin
          CICC1851_compareStage_controlPipe_translated_payload_horizontalDiff = (compareStage_counterOnePixelStream_payload - compareStage_mainOnePixelStream_payload);
        end
      end else begin
        if(when_SuperResolutionPart3_l694) begin
          if(compareStage_controlPipe_payload_horizontalCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_horizontalDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterTwoPixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_horizontalDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainTwoPixelStream_payload);
          end
        end else begin
          if(compareStage_controlPipe_payload_horizontalCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_horizontalDiff = (compareStage_mainThreePixelStream_payload - compareStage_counterThreePixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_horizontalDiff = (compareStage_counterThreePixelStream_payload - compareStage_mainThreePixelStream_payload);
          end
        end
      end
    end
  end

  always @(*) begin
    CICC1851_compareStage_controlPipe_translated_payload_verticalDiff = compareStage_controlPipe_payload_verticalDiff;
    if(compareStage_controlPipe_payload_finalResult) begin
      if(when_SuperResolutionPart3_l647) begin
        CICC1851_compareStage_controlPipe_translated_payload_verticalDiff = 8'h0;
      end else begin
        if(when_SuperResolutionPart3_l649) begin
          if(compareStage_controlPipe_payload_verticalCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_verticalDiff = (compareStage_mainTwoPixelStream_payload - compareStage_mainThreePixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_verticalDiff = (compareStage_mainThreePixelStream_payload - compareStage_mainTwoPixelStream_payload);
          end
        end else begin
          if(when_SuperResolutionPart3_l652) begin
            if(compareStage_controlPipe_payload_verticalCompare) begin
              CICC1851_compareStage_controlPipe_translated_payload_verticalDiff = (compareStage_mainOnePixelStream_payload - compareStage_mainThreePixelStream_payload);
            end else begin
              CICC1851_compareStage_controlPipe_translated_payload_verticalDiff = (compareStage_mainThreePixelStream_payload - compareStage_mainOnePixelStream_payload);
            end
          end else begin
            if(compareStage_controlPipe_payload_verticalCompare) begin
              CICC1851_compareStage_controlPipe_translated_payload_verticalDiff = (compareStage_mainOnePixelStream_payload - compareStage_mainTwoPixelStream_payload);
            end else begin
              CICC1851_compareStage_controlPipe_translated_payload_verticalDiff = (compareStage_mainTwoPixelStream_payload - compareStage_mainOnePixelStream_payload);
            end
          end
        end
      end
    end
  end

  always @(*) begin
    CICC1851_compareStage_controlPipe_translated_payload_inValidMinDiff = compareStage_controlPipe_payload_inValidMinDiff;
    if(when_SuperResolutionPart3_l753) begin
      CICC1851_compareStage_controlPipe_translated_payload_inValidMinDiff = 1'b1;
    end
  end

  assign when_SuperResolutionPart3_l647 = (compareStage_controlPipe_payload_firstRow || compareStage_controlPipe_payload_lastRow);
  assign when_SuperResolutionPart3_l649 = (compareStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l652 = (compareStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l661 = (compareStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l664 = (compareStage_controlPipe_payload_nextPosition == 2'b01);
  assign when_SuperResolutionPart3_l697 = (compareStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l725 = (compareStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l694 = (compareStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l753 = ((((! compareStage_controlPipe_payload_finalResult) && (! compareStage_controlPipe_payload_mainDirectionValid)) && (! compareStage_controlPipe_payload_counterDirectionValid)) && (! compareStage_controlPipe_payload_horizontalDirectionValid));
  assign compareStage_controlPipe_translated_valid = compareStage_controlPipe_valid;
  assign compareStage_controlPipe_ready = compareStage_controlPipe_translated_ready;
  assign compareStage_controlPipe_translated_payload_frameStart = compareStage_controlPipe_payload_frameStart;
  assign compareStage_controlPipe_translated_payload_rowEnd = compareStage_controlPipe_payload_rowEnd;
  assign compareStage_controlPipe_translated_payload_pipeValid = compareStage_controlPipe_payload_pipeValid;
  assign compareStage_controlPipe_translated_payload_firstRow = compareStage_controlPipe_payload_firstRow;
  assign compareStage_controlPipe_translated_payload_lastRow = compareStage_controlPipe_payload_lastRow;
  assign compareStage_controlPipe_translated_payload_finalResult = compareStage_controlPipe_payload_finalResult;
  assign compareStage_controlPipe_translated_payload_mainCompare = compareStage_controlPipe_payload_mainCompare;
  assign compareStage_controlPipe_translated_payload_counterCompare = compareStage_controlPipe_payload_counterCompare;
  assign compareStage_controlPipe_translated_payload_horizontalCompare = compareStage_controlPipe_payload_horizontalCompare;
  assign compareStage_controlPipe_translated_payload_verticalCompare = compareStage_controlPipe_payload_verticalCompare;
  assign compareStage_controlPipe_translated_payload_mainDiff = CICC1851_compareStage_controlPipe_translated_payload_mainDiff;
  assign compareStage_controlPipe_translated_payload_counterDiff = CICC1851_compareStage_controlPipe_translated_payload_counterDiff;
  assign compareStage_controlPipe_translated_payload_horizontalDiff = CICC1851_compareStage_controlPipe_translated_payload_horizontalDiff;
  assign compareStage_controlPipe_translated_payload_verticalDiff = CICC1851_compareStage_controlPipe_translated_payload_verticalDiff;
  assign compareStage_controlPipe_translated_payload_isHorizontalMin = compareStage_controlPipe_payload_isHorizontalMin;
  assign compareStage_controlPipe_translated_payload_minDiff = compareStage_controlPipe_payload_minDiff;
  assign compareStage_controlPipe_translated_payload_currentPosition = compareStage_controlPipe_payload_currentPosition;
  assign compareStage_controlPipe_translated_payload_nextPosition = compareStage_controlPipe_payload_nextPosition;
  assign compareStage_controlPipe_translated_payload_horizontalDirectionValid = compareStage_controlPipe_payload_horizontalDirectionValid;
  assign compareStage_controlPipe_translated_payload_verticalDirectionValid = compareStage_controlPipe_payload_verticalDirectionValid;
  assign compareStage_controlPipe_translated_payload_mainDirectionValid = compareStage_controlPipe_payload_mainDirectionValid;
  assign compareStage_controlPipe_translated_payload_counterDirectionValid = compareStage_controlPipe_payload_counterDirectionValid;
  assign compareStage_controlPipe_translated_payload_inValidMinDiff = CICC1851_compareStage_controlPipe_translated_payload_inValidMinDiff;
  assign compareStage_controlPipe_translated_ready = (! compareStage_controlPipe_translated_rValid);
  assign compareStage_controlPipe_translated_s2mPipe_valid = (compareStage_controlPipe_translated_valid || compareStage_controlPipe_translated_rValid);
  assign compareStage_controlPipe_translated_s2mPipe_payload_frameStart = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_frameStart : compareStage_controlPipe_translated_payload_frameStart);
  assign compareStage_controlPipe_translated_s2mPipe_payload_rowEnd = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_rowEnd : compareStage_controlPipe_translated_payload_rowEnd);
  assign compareStage_controlPipe_translated_s2mPipe_payload_pipeValid = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_pipeValid : compareStage_controlPipe_translated_payload_pipeValid);
  assign compareStage_controlPipe_translated_s2mPipe_payload_firstRow = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_firstRow : compareStage_controlPipe_translated_payload_firstRow);
  assign compareStage_controlPipe_translated_s2mPipe_payload_lastRow = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_lastRow : compareStage_controlPipe_translated_payload_lastRow);
  assign compareStage_controlPipe_translated_s2mPipe_payload_finalResult = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_finalResult : compareStage_controlPipe_translated_payload_finalResult);
  assign compareStage_controlPipe_translated_s2mPipe_payload_mainCompare = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_mainCompare : compareStage_controlPipe_translated_payload_mainCompare);
  assign compareStage_controlPipe_translated_s2mPipe_payload_counterCompare = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_counterCompare : compareStage_controlPipe_translated_payload_counterCompare);
  assign compareStage_controlPipe_translated_s2mPipe_payload_horizontalCompare = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_horizontalCompare : compareStage_controlPipe_translated_payload_horizontalCompare);
  assign compareStage_controlPipe_translated_s2mPipe_payload_verticalCompare = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_verticalCompare : compareStage_controlPipe_translated_payload_verticalCompare);
  assign compareStage_controlPipe_translated_s2mPipe_payload_mainDiff = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_mainDiff : compareStage_controlPipe_translated_payload_mainDiff);
  assign compareStage_controlPipe_translated_s2mPipe_payload_counterDiff = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_counterDiff : compareStage_controlPipe_translated_payload_counterDiff);
  assign compareStage_controlPipe_translated_s2mPipe_payload_horizontalDiff = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_horizontalDiff : compareStage_controlPipe_translated_payload_horizontalDiff);
  assign compareStage_controlPipe_translated_s2mPipe_payload_verticalDiff = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_verticalDiff : compareStage_controlPipe_translated_payload_verticalDiff);
  assign compareStage_controlPipe_translated_s2mPipe_payload_isHorizontalMin = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_isHorizontalMin : compareStage_controlPipe_translated_payload_isHorizontalMin);
  assign compareStage_controlPipe_translated_s2mPipe_payload_minDiff = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_minDiff : compareStage_controlPipe_translated_payload_minDiff);
  assign compareStage_controlPipe_translated_s2mPipe_payload_currentPosition = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_currentPosition : compareStage_controlPipe_translated_payload_currentPosition);
  assign compareStage_controlPipe_translated_s2mPipe_payload_nextPosition = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_nextPosition : compareStage_controlPipe_translated_payload_nextPosition);
  assign compareStage_controlPipe_translated_s2mPipe_payload_horizontalDirectionValid = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_horizontalDirectionValid : compareStage_controlPipe_translated_payload_horizontalDirectionValid);
  assign compareStage_controlPipe_translated_s2mPipe_payload_verticalDirectionValid = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_verticalDirectionValid : compareStage_controlPipe_translated_payload_verticalDirectionValid);
  assign compareStage_controlPipe_translated_s2mPipe_payload_mainDirectionValid = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_mainDirectionValid : compareStage_controlPipe_translated_payload_mainDirectionValid);
  assign compareStage_controlPipe_translated_s2mPipe_payload_counterDirectionValid = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_counterDirectionValid : compareStage_controlPipe_translated_payload_counterDirectionValid);
  assign compareStage_controlPipe_translated_s2mPipe_payload_inValidMinDiff = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_inValidMinDiff : compareStage_controlPipe_translated_payload_inValidMinDiff);
  always @(*) begin
    compareStage_controlPipe_translated_s2mPipe_ready = diffStage_controlPipe_ready;
    if(when_Stream_l368_53) begin
      compareStage_controlPipe_translated_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_53 = (! diffStage_controlPipe_valid);
  assign diffStage_controlPipe_valid = compareStage_controlPipe_translated_s2mPipe_rValid;
  assign diffStage_controlPipe_payload_frameStart = compareStage_controlPipe_translated_s2mPipe_rData_frameStart;
  assign diffStage_controlPipe_payload_rowEnd = compareStage_controlPipe_translated_s2mPipe_rData_rowEnd;
  assign diffStage_controlPipe_payload_pipeValid = compareStage_controlPipe_translated_s2mPipe_rData_pipeValid;
  assign diffStage_controlPipe_payload_firstRow = compareStage_controlPipe_translated_s2mPipe_rData_firstRow;
  assign diffStage_controlPipe_payload_lastRow = compareStage_controlPipe_translated_s2mPipe_rData_lastRow;
  assign diffStage_controlPipe_payload_finalResult = compareStage_controlPipe_translated_s2mPipe_rData_finalResult;
  assign diffStage_controlPipe_payload_mainCompare = compareStage_controlPipe_translated_s2mPipe_rData_mainCompare;
  assign diffStage_controlPipe_payload_counterCompare = compareStage_controlPipe_translated_s2mPipe_rData_counterCompare;
  assign diffStage_controlPipe_payload_horizontalCompare = compareStage_controlPipe_translated_s2mPipe_rData_horizontalCompare;
  assign diffStage_controlPipe_payload_verticalCompare = compareStage_controlPipe_translated_s2mPipe_rData_verticalCompare;
  assign diffStage_controlPipe_payload_mainDiff = compareStage_controlPipe_translated_s2mPipe_rData_mainDiff;
  assign diffStage_controlPipe_payload_counterDiff = compareStage_controlPipe_translated_s2mPipe_rData_counterDiff;
  assign diffStage_controlPipe_payload_horizontalDiff = compareStage_controlPipe_translated_s2mPipe_rData_horizontalDiff;
  assign diffStage_controlPipe_payload_verticalDiff = compareStage_controlPipe_translated_s2mPipe_rData_verticalDiff;
  assign diffStage_controlPipe_payload_isHorizontalMin = compareStage_controlPipe_translated_s2mPipe_rData_isHorizontalMin;
  assign diffStage_controlPipe_payload_minDiff = compareStage_controlPipe_translated_s2mPipe_rData_minDiff;
  assign diffStage_controlPipe_payload_currentPosition = compareStage_controlPipe_translated_s2mPipe_rData_currentPosition;
  assign diffStage_controlPipe_payload_nextPosition = compareStage_controlPipe_translated_s2mPipe_rData_nextPosition;
  assign diffStage_controlPipe_payload_horizontalDirectionValid = compareStage_controlPipe_translated_s2mPipe_rData_horizontalDirectionValid;
  assign diffStage_controlPipe_payload_verticalDirectionValid = compareStage_controlPipe_translated_s2mPipe_rData_verticalDirectionValid;
  assign diffStage_controlPipe_payload_mainDirectionValid = compareStage_controlPipe_translated_s2mPipe_rData_mainDirectionValid;
  assign diffStage_controlPipe_payload_counterDirectionValid = compareStage_controlPipe_translated_s2mPipe_rData_counterDirectionValid;
  assign diffStage_controlPipe_payload_inValidMinDiff = compareStage_controlPipe_translated_s2mPipe_rData_inValidMinDiff;
  assign diffStage_mainOnePixelStream_ready = (! diffStage_mainOnePixelStream_rValid);
  assign diffStage_mainOnePixelStream_s2mPipe_valid = (diffStage_mainOnePixelStream_valid || diffStage_mainOnePixelStream_rValid);
  assign diffStage_mainOnePixelStream_s2mPipe_payload = (diffStage_mainOnePixelStream_rValid ? diffStage_mainOnePixelStream_rData : diffStage_mainOnePixelStream_payload);
  always @(*) begin
    diffStage_mainOnePixelStream_s2mPipe_ready = resultStage_mainOnePixelStream_ready;
    if(when_Stream_l368_54) begin
      diffStage_mainOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_54 = (! resultStage_mainOnePixelStream_valid);
  assign resultStage_mainOnePixelStream_valid = diffStage_mainOnePixelStream_s2mPipe_rValid;
  assign resultStage_mainOnePixelStream_payload = diffStage_mainOnePixelStream_s2mPipe_rData;
  assign diffStage_counterOnePixelStream_ready = (! diffStage_counterOnePixelStream_rValid);
  assign diffStage_counterOnePixelStream_s2mPipe_valid = (diffStage_counterOnePixelStream_valid || diffStage_counterOnePixelStream_rValid);
  assign diffStage_counterOnePixelStream_s2mPipe_payload = (diffStage_counterOnePixelStream_rValid ? diffStage_counterOnePixelStream_rData : diffStage_counterOnePixelStream_payload);
  always @(*) begin
    diffStage_counterOnePixelStream_s2mPipe_ready = resultStage_counterOnePixelStream_ready;
    if(when_Stream_l368_55) begin
      diffStage_counterOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_55 = (! resultStage_counterOnePixelStream_valid);
  assign resultStage_counterOnePixelStream_valid = diffStage_counterOnePixelStream_s2mPipe_rValid;
  assign resultStage_counterOnePixelStream_payload = diffStage_counterOnePixelStream_s2mPipe_rData;
  assign diffStage_mainTwoPixelStream_ready = (! diffStage_mainTwoPixelStream_rValid);
  assign diffStage_mainTwoPixelStream_s2mPipe_valid = (diffStage_mainTwoPixelStream_valid || diffStage_mainTwoPixelStream_rValid);
  assign diffStage_mainTwoPixelStream_s2mPipe_payload = (diffStage_mainTwoPixelStream_rValid ? diffStage_mainTwoPixelStream_rData : diffStage_mainTwoPixelStream_payload);
  always @(*) begin
    diffStage_mainTwoPixelStream_s2mPipe_ready = resultStage_mainTwoPixelStream_ready;
    if(when_Stream_l368_56) begin
      diffStage_mainTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_56 = (! resultStage_mainTwoPixelStream_valid);
  assign resultStage_mainTwoPixelStream_valid = diffStage_mainTwoPixelStream_s2mPipe_rValid;
  assign resultStage_mainTwoPixelStream_payload = diffStage_mainTwoPixelStream_s2mPipe_rData;
  assign diffStage_counterTwoPixelStream_ready = (! diffStage_counterTwoPixelStream_rValid);
  assign diffStage_counterTwoPixelStream_s2mPipe_valid = (diffStage_counterTwoPixelStream_valid || diffStage_counterTwoPixelStream_rValid);
  assign diffStage_counterTwoPixelStream_s2mPipe_payload = (diffStage_counterTwoPixelStream_rValid ? diffStage_counterTwoPixelStream_rData : diffStage_counterTwoPixelStream_payload);
  always @(*) begin
    diffStage_counterTwoPixelStream_s2mPipe_ready = resultStage_counterTwoPixelStream_ready;
    if(when_Stream_l368_57) begin
      diffStage_counterTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_57 = (! resultStage_counterTwoPixelStream_valid);
  assign resultStage_counterTwoPixelStream_valid = diffStage_counterTwoPixelStream_s2mPipe_rValid;
  assign resultStage_counterTwoPixelStream_payload = diffStage_counterTwoPixelStream_s2mPipe_rData;
  assign diffStage_mainThreePixelStream_ready = (! diffStage_mainThreePixelStream_rValid);
  assign diffStage_mainThreePixelStream_s2mPipe_valid = (diffStage_mainThreePixelStream_valid || diffStage_mainThreePixelStream_rValid);
  assign diffStage_mainThreePixelStream_s2mPipe_payload = (diffStage_mainThreePixelStream_rValid ? diffStage_mainThreePixelStream_rData : diffStage_mainThreePixelStream_payload);
  always @(*) begin
    diffStage_mainThreePixelStream_s2mPipe_ready = resultStage_mainThreePixelStream_ready;
    if(when_Stream_l368_58) begin
      diffStage_mainThreePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_58 = (! resultStage_mainThreePixelStream_valid);
  assign resultStage_mainThreePixelStream_valid = diffStage_mainThreePixelStream_s2mPipe_rValid;
  assign resultStage_mainThreePixelStream_payload = diffStage_mainThreePixelStream_s2mPipe_rData;
  assign diffStage_counterThreePixelStream_ready = (! diffStage_counterThreePixelStream_rValid);
  assign diffStage_counterThreePixelStream_s2mPipe_valid = (diffStage_counterThreePixelStream_valid || diffStage_counterThreePixelStream_rValid);
  assign diffStage_counterThreePixelStream_s2mPipe_payload = (diffStage_counterThreePixelStream_rValid ? diffStage_counterThreePixelStream_rData : diffStage_counterThreePixelStream_payload);
  always @(*) begin
    diffStage_counterThreePixelStream_s2mPipe_ready = resultStage_counterThreePixelStream_ready;
    if(when_Stream_l368_59) begin
      diffStage_counterThreePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_59 = (! resultStage_counterThreePixelStream_valid);
  assign resultStage_counterThreePixelStream_valid = diffStage_counterThreePixelStream_s2mPipe_rValid;
  assign resultStage_counterThreePixelStream_payload = diffStage_counterThreePixelStream_s2mPipe_rData;
  assign diffStage_mainOneValidStream_ready = (! diffStage_mainOneValidStream_rValid);
  assign diffStage_mainOneValidStream_s2mPipe_valid = (diffStage_mainOneValidStream_valid || diffStage_mainOneValidStream_rValid);
  assign diffStage_mainOneValidStream_s2mPipe_payload = (diffStage_mainOneValidStream_rValid ? diffStage_mainOneValidStream_rData : diffStage_mainOneValidStream_payload);
  always @(*) begin
    diffStage_mainOneValidStream_s2mPipe_ready = resultStage_mainOneValidStream_ready;
    if(when_Stream_l368_60) begin
      diffStage_mainOneValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_60 = (! resultStage_mainOneValidStream_valid);
  assign resultStage_mainOneValidStream_valid = diffStage_mainOneValidStream_s2mPipe_rValid;
  assign resultStage_mainOneValidStream_payload = diffStage_mainOneValidStream_s2mPipe_rData;
  assign diffStage_counterOneValidStream_ready = (! diffStage_counterOneValidStream_rValid);
  assign diffStage_counterOneValidStream_s2mPipe_valid = (diffStage_counterOneValidStream_valid || diffStage_counterOneValidStream_rValid);
  assign diffStage_counterOneValidStream_s2mPipe_payload = (diffStage_counterOneValidStream_rValid ? diffStage_counterOneValidStream_rData : diffStage_counterOneValidStream_payload);
  always @(*) begin
    diffStage_counterOneValidStream_s2mPipe_ready = resultStage_counterOneValidStream_ready;
    if(when_Stream_l368_61) begin
      diffStage_counterOneValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_61 = (! resultStage_counterOneValidStream_valid);
  assign resultStage_counterOneValidStream_valid = diffStage_counterOneValidStream_s2mPipe_rValid;
  assign resultStage_counterOneValidStream_payload = diffStage_counterOneValidStream_s2mPipe_rData;
  assign diffStage_mainTwoValidStream_ready = (! diffStage_mainTwoValidStream_rValid);
  assign diffStage_mainTwoValidStream_s2mPipe_valid = (diffStage_mainTwoValidStream_valid || diffStage_mainTwoValidStream_rValid);
  assign diffStage_mainTwoValidStream_s2mPipe_payload = (diffStage_mainTwoValidStream_rValid ? diffStage_mainTwoValidStream_rData : diffStage_mainTwoValidStream_payload);
  always @(*) begin
    diffStage_mainTwoValidStream_s2mPipe_ready = resultStage_mainTwoValidStream_ready;
    if(when_Stream_l368_62) begin
      diffStage_mainTwoValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_62 = (! resultStage_mainTwoValidStream_valid);
  assign resultStage_mainTwoValidStream_valid = diffStage_mainTwoValidStream_s2mPipe_rValid;
  assign resultStage_mainTwoValidStream_payload = diffStage_mainTwoValidStream_s2mPipe_rData;
  assign diffStage_counterTwoValidStream_ready = (! diffStage_counterTwoValidStream_rValid);
  assign diffStage_counterTwoValidStream_s2mPipe_valid = (diffStage_counterTwoValidStream_valid || diffStage_counterTwoValidStream_rValid);
  assign diffStage_counterTwoValidStream_s2mPipe_payload = (diffStage_counterTwoValidStream_rValid ? diffStage_counterTwoValidStream_rData : diffStage_counterTwoValidStream_payload);
  always @(*) begin
    diffStage_counterTwoValidStream_s2mPipe_ready = resultStage_counterTwoValidStream_ready;
    if(when_Stream_l368_63) begin
      diffStage_counterTwoValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_63 = (! resultStage_counterTwoValidStream_valid);
  assign resultStage_counterTwoValidStream_valid = diffStage_counterTwoValidStream_s2mPipe_rValid;
  assign resultStage_counterTwoValidStream_payload = diffStage_counterTwoValidStream_s2mPipe_rData;
  assign diffStage_mainThreeValidStream_ready = (! diffStage_mainThreeValidStream_rValid);
  assign diffStage_mainThreeValidStream_s2mPipe_valid = (diffStage_mainThreeValidStream_valid || diffStage_mainThreeValidStream_rValid);
  assign diffStage_mainThreeValidStream_s2mPipe_payload = (diffStage_mainThreeValidStream_rValid ? diffStage_mainThreeValidStream_rData : diffStage_mainThreeValidStream_payload);
  always @(*) begin
    diffStage_mainThreeValidStream_s2mPipe_ready = resultStage_mainThreeValidStream_ready;
    if(when_Stream_l368_64) begin
      diffStage_mainThreeValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_64 = (! resultStage_mainThreeValidStream_valid);
  assign resultStage_mainThreeValidStream_valid = diffStage_mainThreeValidStream_s2mPipe_rValid;
  assign resultStage_mainThreeValidStream_payload = diffStage_mainThreeValidStream_s2mPipe_rData;
  assign diffStage_counterThreeValidStream_ready = (! diffStage_counterThreeValidStream_rValid);
  assign diffStage_counterThreeValidStream_s2mPipe_valid = (diffStage_counterThreeValidStream_valid || diffStage_counterThreeValidStream_rValid);
  assign diffStage_counterThreeValidStream_s2mPipe_payload = (diffStage_counterThreeValidStream_rValid ? diffStage_counterThreeValidStream_rData : diffStage_counterThreeValidStream_payload);
  always @(*) begin
    diffStage_counterThreeValidStream_s2mPipe_ready = resultStage_counterThreeValidStream_ready;
    if(when_Stream_l368_65) begin
      diffStage_counterThreeValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_65 = (! resultStage_counterThreeValidStream_valid);
  assign resultStage_counterThreeValidStream_valid = diffStage_counterThreeValidStream_s2mPipe_rValid;
  assign resultStage_counterThreeValidStream_payload = diffStage_counterThreeValidStream_s2mPipe_rData;
  assign diffStage_controlPipe_ready = diffStage_controlPipe_fork_io_input_ready;
  always @(*) begin
    CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin = diffStage_controlPipe_payload_isHorizontalMin;
    if(when_SuperResolutionPart3_l783) begin
      if(when_SuperResolutionPart3_l784) begin
        if(when_SuperResolutionPart3_l785) begin
          CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin = 1'b1;
        end else begin
          if(when_SuperResolutionPart3_l788) begin
            CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin = 1'b0;
          end else begin
            CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin = 1'b0;
          end
        end
      end else begin
        if(when_SuperResolutionPart3_l795) begin
          if(when_SuperResolutionPart3_l796) begin
            CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin = 1'b0;
          end else begin
            CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin = 1'b0;
          end
        end else begin
          if(when_SuperResolutionPart3_l803) begin
            if(when_SuperResolutionPart3_l804) begin
              CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin = 1'b1;
            end else begin
              CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin = 1'b0;
            end
          end else begin
            if(when_SuperResolutionPart3_l811) begin
              if(when_SuperResolutionPart3_l812) begin
                CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin = 1'b1;
              end else begin
                CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l819) begin
                CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin = 1'b0;
              end else begin
                if(when_SuperResolutionPart3_l822) begin
                  CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin = 1'b1;
                end else begin
                  if(when_SuperResolutionPart3_l825) begin
                    CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin = 1'b0;
                  end
                end
              end
            end
          end
        end
      end
    end
  end

  always @(*) begin
    CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff = diffStage_controlPipe_payload_minDiff;
    if(when_SuperResolutionPart3_l783) begin
      if(when_SuperResolutionPart3_l784) begin
        if(when_SuperResolutionPart3_l785) begin
          CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff = diffStage_controlPipe_payload_horizontalDiff;
        end else begin
          if(when_SuperResolutionPart3_l788) begin
            CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff = diffStage_controlPipe_payload_mainDiff;
          end else begin
            CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff = diffStage_controlPipe_payload_counterDiff;
          end
        end
      end else begin
        if(when_SuperResolutionPart3_l795) begin
          if(when_SuperResolutionPart3_l796) begin
            CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff = diffStage_controlPipe_payload_mainDiff;
          end else begin
            CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff = diffStage_controlPipe_payload_counterDiff;
          end
        end else begin
          if(when_SuperResolutionPart3_l803) begin
            if(when_SuperResolutionPart3_l804) begin
              CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff = diffStage_controlPipe_payload_horizontalDiff;
            end else begin
              CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff = diffStage_controlPipe_payload_counterDiff;
            end
          end else begin
            if(when_SuperResolutionPart3_l811) begin
              if(when_SuperResolutionPart3_l812) begin
                CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff = diffStage_controlPipe_payload_horizontalDiff;
              end else begin
                CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff = diffStage_controlPipe_payload_mainDiff;
              end
            end else begin
              if(when_SuperResolutionPart3_l819) begin
                CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff = diffStage_controlPipe_payload_counterDiff;
              end else begin
                if(when_SuperResolutionPart3_l822) begin
                  CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff = diffStage_controlPipe_payload_horizontalDiff;
                end else begin
                  if(when_SuperResolutionPart3_l825) begin
                    CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff = diffStage_controlPipe_payload_mainDiff;
                  end
                end
              end
            end
          end
        end
      end
    end
  end

  assign when_SuperResolutionPart3_l783 = (! diffStage_controlPipe_payload_finalResult);
  assign when_SuperResolutionPart3_l784 = ((diffStage_controlPipe_payload_horizontalDirectionValid && diffStage_controlPipe_payload_mainDirectionValid) && diffStage_controlPipe_payload_counterDirectionValid);
  assign when_SuperResolutionPart3_l785 = ((diffStage_controlPipe_payload_horizontalDiff <= diffStage_controlPipe_payload_mainDiff) && (diffStage_controlPipe_payload_horizontalDiff <= diffStage_controlPipe_payload_counterDiff));
  assign when_SuperResolutionPart3_l788 = ((diffStage_controlPipe_payload_mainDiff < diffStage_controlPipe_payload_horizontalDiff) && (diffStage_controlPipe_payload_mainDiff <= diffStage_controlPipe_payload_counterDiff));
  assign when_SuperResolutionPart3_l796 = (diffStage_controlPipe_payload_mainDiff <= diffStage_controlPipe_payload_counterDiff);
  assign when_SuperResolutionPart3_l804 = (diffStage_controlPipe_payload_horizontalDiff <= diffStage_controlPipe_payload_counterDiff);
  assign when_SuperResolutionPart3_l812 = (diffStage_controlPipe_payload_horizontalDiff <= diffStage_controlPipe_payload_mainDiff);
  assign when_SuperResolutionPart3_l795 = (((! diffStage_controlPipe_payload_horizontalDirectionValid) && diffStage_controlPipe_payload_mainDirectionValid) && diffStage_controlPipe_payload_counterDirectionValid);
  assign when_SuperResolutionPart3_l803 = ((diffStage_controlPipe_payload_horizontalDirectionValid && (! diffStage_controlPipe_payload_mainDirectionValid)) && diffStage_controlPipe_payload_counterDirectionValid);
  assign when_SuperResolutionPart3_l811 = ((diffStage_controlPipe_payload_horizontalDirectionValid && diffStage_controlPipe_payload_mainDirectionValid) && (! diffStage_controlPipe_payload_counterDirectionValid));
  assign when_SuperResolutionPart3_l819 = (((! diffStage_controlPipe_payload_horizontalDirectionValid) && (! diffStage_controlPipe_payload_mainDirectionValid)) && diffStage_controlPipe_payload_counterDirectionValid);
  assign when_SuperResolutionPart3_l822 = ((diffStage_controlPipe_payload_horizontalDirectionValid && (! diffStage_controlPipe_payload_mainDirectionValid)) && (! diffStage_controlPipe_payload_counterDirectionValid));
  assign when_SuperResolutionPart3_l825 = (((! diffStage_controlPipe_payload_horizontalDirectionValid) && diffStage_controlPipe_payload_mainDirectionValid) && (! diffStage_controlPipe_payload_counterDirectionValid));
  assign resultStage_controlPipeBeforePipe_valid = diffStage_controlPipe_fork_io_outputs_0_valid;
  assign resultStage_controlPipeBeforePipe_payload_frameStart = diffStage_controlPipe_payload_frameStart;
  assign resultStage_controlPipeBeforePipe_payload_rowEnd = diffStage_controlPipe_payload_rowEnd;
  assign resultStage_controlPipeBeforePipe_payload_pipeValid = diffStage_controlPipe_payload_pipeValid;
  assign resultStage_controlPipeBeforePipe_payload_firstRow = diffStage_controlPipe_payload_firstRow;
  assign resultStage_controlPipeBeforePipe_payload_lastRow = diffStage_controlPipe_payload_lastRow;
  assign resultStage_controlPipeBeforePipe_payload_finalResult = diffStage_controlPipe_payload_finalResult;
  assign resultStage_controlPipeBeforePipe_payload_mainCompare = diffStage_controlPipe_payload_mainCompare;
  assign resultStage_controlPipeBeforePipe_payload_counterCompare = diffStage_controlPipe_payload_counterCompare;
  assign resultStage_controlPipeBeforePipe_payload_horizontalCompare = diffStage_controlPipe_payload_horizontalCompare;
  assign resultStage_controlPipeBeforePipe_payload_verticalCompare = diffStage_controlPipe_payload_verticalCompare;
  assign resultStage_controlPipeBeforePipe_payload_mainDiff = diffStage_controlPipe_payload_mainDiff;
  assign resultStage_controlPipeBeforePipe_payload_counterDiff = diffStage_controlPipe_payload_counterDiff;
  assign resultStage_controlPipeBeforePipe_payload_horizontalDiff = diffStage_controlPipe_payload_horizontalDiff;
  assign resultStage_controlPipeBeforePipe_payload_verticalDiff = diffStage_controlPipe_payload_verticalDiff;
  assign resultStage_controlPipeBeforePipe_payload_isHorizontalMin = CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin;
  assign resultStage_controlPipeBeforePipe_payload_minDiff = CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff;
  assign resultStage_controlPipeBeforePipe_payload_currentPosition = diffStage_controlPipe_payload_currentPosition;
  assign resultStage_controlPipeBeforePipe_payload_nextPosition = diffStage_controlPipe_payload_nextPosition;
  assign resultStage_controlPipeBeforePipe_payload_horizontalDirectionValid = diffStage_controlPipe_payload_horizontalDirectionValid;
  assign resultStage_controlPipeBeforePipe_payload_verticalDirectionValid = diffStage_controlPipe_payload_verticalDirectionValid;
  assign resultStage_controlPipeBeforePipe_payload_mainDirectionValid = diffStage_controlPipe_payload_mainDirectionValid;
  assign resultStage_controlPipeBeforePipe_payload_counterDirectionValid = diffStage_controlPipe_payload_counterDirectionValid;
  assign resultStage_controlPipeBeforePipe_payload_inValidMinDiff = diffStage_controlPipe_payload_inValidMinDiff;
  assign resultStage_controlPipeBeforePipe_ready = (! resultStage_controlPipeBeforePipe_rValid);
  assign resultStage_controlPipeBeforePipe_s2mPipe_valid = (resultStage_controlPipeBeforePipe_valid || resultStage_controlPipeBeforePipe_rValid);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_frameStart = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_frameStart : resultStage_controlPipeBeforePipe_payload_frameStart);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_rowEnd = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_rowEnd : resultStage_controlPipeBeforePipe_payload_rowEnd);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_pipeValid = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_pipeValid : resultStage_controlPipeBeforePipe_payload_pipeValid);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_firstRow = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_firstRow : resultStage_controlPipeBeforePipe_payload_firstRow);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_lastRow = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_lastRow : resultStage_controlPipeBeforePipe_payload_lastRow);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_finalResult = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_finalResult : resultStage_controlPipeBeforePipe_payload_finalResult);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_mainCompare = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_mainCompare : resultStage_controlPipeBeforePipe_payload_mainCompare);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_counterCompare = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_counterCompare : resultStage_controlPipeBeforePipe_payload_counterCompare);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_horizontalCompare = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_horizontalCompare : resultStage_controlPipeBeforePipe_payload_horizontalCompare);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_verticalCompare = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_verticalCompare : resultStage_controlPipeBeforePipe_payload_verticalCompare);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_mainDiff = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_mainDiff : resultStage_controlPipeBeforePipe_payload_mainDiff);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_counterDiff = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_counterDiff : resultStage_controlPipeBeforePipe_payload_counterDiff);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_horizontalDiff = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_horizontalDiff : resultStage_controlPipeBeforePipe_payload_horizontalDiff);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_verticalDiff = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_verticalDiff : resultStage_controlPipeBeforePipe_payload_verticalDiff);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_isHorizontalMin = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_isHorizontalMin : resultStage_controlPipeBeforePipe_payload_isHorizontalMin);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_minDiff = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_minDiff : resultStage_controlPipeBeforePipe_payload_minDiff);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_currentPosition = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_currentPosition : resultStage_controlPipeBeforePipe_payload_currentPosition);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_nextPosition = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_nextPosition : resultStage_controlPipeBeforePipe_payload_nextPosition);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_horizontalDirectionValid = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_horizontalDirectionValid : resultStage_controlPipeBeforePipe_payload_horizontalDirectionValid);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_verticalDirectionValid = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_verticalDirectionValid : resultStage_controlPipeBeforePipe_payload_verticalDirectionValid);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_mainDirectionValid = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_mainDirectionValid : resultStage_controlPipeBeforePipe_payload_mainDirectionValid);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_counterDirectionValid = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_counterDirectionValid : resultStage_controlPipeBeforePipe_payload_counterDirectionValid);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_inValidMinDiff = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_inValidMinDiff : resultStage_controlPipeBeforePipe_payload_inValidMinDiff);
  always @(*) begin
    resultStage_controlPipeBeforePipe_s2mPipe_ready = resultStage_controlPipe_ready;
    if(when_Stream_l368_66) begin
      resultStage_controlPipeBeforePipe_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_66 = (! resultStage_controlPipe_valid);
  assign resultStage_controlPipe_valid = resultStage_controlPipeBeforePipe_s2mPipe_rValid;
  assign resultStage_controlPipe_payload_frameStart = resultStage_controlPipeBeforePipe_s2mPipe_rData_frameStart;
  assign resultStage_controlPipe_payload_rowEnd = resultStage_controlPipeBeforePipe_s2mPipe_rData_rowEnd;
  assign resultStage_controlPipe_payload_pipeValid = resultStage_controlPipeBeforePipe_s2mPipe_rData_pipeValid;
  assign resultStage_controlPipe_payload_firstRow = resultStage_controlPipeBeforePipe_s2mPipe_rData_firstRow;
  assign resultStage_controlPipe_payload_lastRow = resultStage_controlPipeBeforePipe_s2mPipe_rData_lastRow;
  assign resultStage_controlPipe_payload_finalResult = resultStage_controlPipeBeforePipe_s2mPipe_rData_finalResult;
  assign resultStage_controlPipe_payload_mainCompare = resultStage_controlPipeBeforePipe_s2mPipe_rData_mainCompare;
  assign resultStage_controlPipe_payload_counterCompare = resultStage_controlPipeBeforePipe_s2mPipe_rData_counterCompare;
  assign resultStage_controlPipe_payload_horizontalCompare = resultStage_controlPipeBeforePipe_s2mPipe_rData_horizontalCompare;
  assign resultStage_controlPipe_payload_verticalCompare = resultStage_controlPipeBeforePipe_s2mPipe_rData_verticalCompare;
  assign resultStage_controlPipe_payload_mainDiff = resultStage_controlPipeBeforePipe_s2mPipe_rData_mainDiff;
  assign resultStage_controlPipe_payload_counterDiff = resultStage_controlPipeBeforePipe_s2mPipe_rData_counterDiff;
  assign resultStage_controlPipe_payload_horizontalDiff = resultStage_controlPipeBeforePipe_s2mPipe_rData_horizontalDiff;
  assign resultStage_controlPipe_payload_verticalDiff = resultStage_controlPipeBeforePipe_s2mPipe_rData_verticalDiff;
  assign resultStage_controlPipe_payload_isHorizontalMin = resultStage_controlPipeBeforePipe_s2mPipe_rData_isHorizontalMin;
  assign resultStage_controlPipe_payload_minDiff = resultStage_controlPipeBeforePipe_s2mPipe_rData_minDiff;
  assign resultStage_controlPipe_payload_currentPosition = resultStage_controlPipeBeforePipe_s2mPipe_rData_currentPosition;
  assign resultStage_controlPipe_payload_nextPosition = resultStage_controlPipeBeforePipe_s2mPipe_rData_nextPosition;
  assign resultStage_controlPipe_payload_horizontalDirectionValid = resultStage_controlPipeBeforePipe_s2mPipe_rData_horizontalDirectionValid;
  assign resultStage_controlPipe_payload_verticalDirectionValid = resultStage_controlPipeBeforePipe_s2mPipe_rData_verticalDirectionValid;
  assign resultStage_controlPipe_payload_mainDirectionValid = resultStage_controlPipeBeforePipe_s2mPipe_rData_mainDirectionValid;
  assign resultStage_controlPipe_payload_counterDirectionValid = resultStage_controlPipeBeforePipe_s2mPipe_rData_counterDirectionValid;
  assign resultStage_controlPipe_payload_inValidMinDiff = resultStage_controlPipeBeforePipe_s2mPipe_rData_inValidMinDiff;
  assign resultStage_pixelStream_valid = diffStage_controlPipe_fork_io_outputs_1_valid;
  always @(*) begin
    resultStage_pixelStream_payload = 8'h0;
    if(diffStage_controlPipe_payload_finalResult) begin
      if(when_SuperResolutionPart3_l840) begin
        resultStage_pixelStream_payload = diffStage_mainOnePixelStream_payload;
      end else begin
        if(when_SuperResolutionPart3_l841) begin
          resultStage_pixelStream_payload = diffStage_mainTwoPixelStream_payload;
        end else begin
          if(when_SuperResolutionPart3_l842) begin
            resultStage_pixelStream_payload = diffStage_mainThreePixelStream_payload;
          end else begin
            if(diffStage_controlPipe_payload_verticalDirectionValid) begin
              if(inValidMinDiff) begin
                if(when_SuperResolutionPart3_l846) begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload[7:0];
                end else begin
                  if(when_SuperResolutionPart3_l847) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_2[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_4[7:0];
                  end
                end
              end else begin
                if(when_SuperResolutionPart3_l850) begin
                  resultStage_pixelStream_payload = candidatePixel;
                end else begin
                  if(when_SuperResolutionPart3_l851) begin
                    if(isHorizontalDirection) begin
                      resultStage_pixelStream_payload = candidatePixel;
                    end else begin
                      if(when_SuperResolutionPart3_l854) begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_6[7:0];
                      end else begin
                        if(when_SuperResolutionPart3_l855) begin
                          resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_8[7:0];
                        end else begin
                          resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_10[7:0];
                        end
                      end
                    end
                  end else begin
                    if(when_SuperResolutionPart3_l860) begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_12[7:0];
                    end else begin
                      if(when_SuperResolutionPart3_l861) begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_14[7:0];
                      end else begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_16[7:0];
                      end
                    end
                  end
                end
              end
            end else begin
              resultStage_pixelStream_payload = candidatePixel;
            end
          end
        end
      end
    end else begin
      if(when_SuperResolutionPart3_l869) begin
        if(when_SuperResolutionPart3_l870) begin
          if(when_SuperResolutionPart3_l871) begin
            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_18[7:0];
          end else begin
            if(when_SuperResolutionPart3_l872) begin
              resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_20[7:0];
            end else begin
              resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_22[7:0];
            end
          end
        end else begin
          if(when_SuperResolutionPart3_l874) begin
            if(when_SuperResolutionPart3_l875) begin
              if(when_SuperResolutionPart3_l876) begin
                if(diffStage_controlPipe_payload_firstRow) begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_24[7:0];
                end else begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_26[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_28[7:0];
                  end
                end
              end else begin
                if(diffStage_controlPipe_payload_lastRow) begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_30[7:0];
                end else begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_32[7:0];
                end
              end
            end else begin
              if(when_SuperResolutionPart3_l884) begin
                if(when_SuperResolutionPart3_l885) begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_34[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_36[7:0];
                  end
                end else begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_38[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_40[7:0];
                  end
                end
              end else begin
                if(when_SuperResolutionPart3_l893) begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_42[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_44[7:0];
                  end
                end else begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_46[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_48[7:0];
                  end
                end
              end
            end
          end else begin
            if(when_SuperResolutionPart3_l902) begin
              if(when_SuperResolutionPart3_l903) begin
                if(diffStage_controlPipe_payload_firstRow) begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_50[7:0];
                end else begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_52[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_54[7:0];
                  end
                end
              end else begin
                if(diffStage_controlPipe_payload_lastRow) begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_56[7:0];
                end else begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_58[7:0];
                end
              end
            end else begin
              if(when_SuperResolutionPart3_l911) begin
                if(when_SuperResolutionPart3_l912) begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_60[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_62[7:0];
                  end
                end else begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_64[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_66[7:0];
                  end
                end
              end else begin
                if(when_SuperResolutionPart3_l920) begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_68[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_70[7:0];
                  end
                end else begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_72[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_74[7:0];
                  end
                end
              end
            end
          end
        end
      end else begin
        if(when_SuperResolutionPart3_l929) begin
          if(when_SuperResolutionPart3_l930) begin
            if(when_SuperResolutionPart3_l931) begin
              if(when_SuperResolutionPart3_l932) begin
                if(diffStage_controlPipe_payload_firstRow) begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_76[7:0];
                end else begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_78[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_80[7:0];
                  end
                end
              end else begin
                if(diffStage_controlPipe_payload_lastRow) begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_82[7:0];
                end else begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_84[7:0];
                end
              end
            end else begin
              if(when_SuperResolutionPart3_l940) begin
                if(when_SuperResolutionPart3_l941) begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_86[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_88[7:0];
                  end
                end else begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_90[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_92[7:0];
                  end
                end
              end else begin
                if(when_SuperResolutionPart3_l949) begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_94[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_96[7:0];
                  end
                end else begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_98[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_100[7:0];
                  end
                end
              end
            end
          end else begin
            if(when_SuperResolutionPart3_l958) begin
              if(when_SuperResolutionPart3_l959) begin
                if(diffStage_controlPipe_payload_firstRow) begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_102[7:0];
                end else begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_104[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_106[7:0];
                  end
                end
              end else begin
                if(diffStage_controlPipe_payload_lastRow) begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_108[7:0];
                end else begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_110[7:0];
                end
              end
            end else begin
              if(when_SuperResolutionPart3_l967) begin
                if(when_SuperResolutionPart3_l968) begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_112[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_114[7:0];
                  end
                end else begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_116[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_118[7:0];
                  end
                end
              end else begin
                if(when_SuperResolutionPart3_l976) begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_120[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_122[7:0];
                  end
                end else begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_124[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_126[7:0];
                  end
                end
              end
            end
          end
        end else begin
          if(when_SuperResolutionPart3_l985) begin
            if(when_SuperResolutionPart3_l986) begin
              if(when_SuperResolutionPart3_l987) begin
                resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_128[7:0];
              end else begin
                if(when_SuperResolutionPart3_l988) begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_130[7:0];
                end else begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_132[7:0];
                end
              end
            end else begin
              if(when_SuperResolutionPart3_l991) begin
                if(when_SuperResolutionPart3_l992) begin
                  if(diffStage_controlPipe_payload_firstRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_134[7:0];
                  end else begin
                    if(diffStage_controlPipe_payload_lastRow) begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_136[7:0];
                    end else begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_138[7:0];
                    end
                  end
                end else begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_140[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_142[7:0];
                  end
                end
              end else begin
                if(when_SuperResolutionPart3_l1000) begin
                  if(when_SuperResolutionPart3_l1001) begin
                    if(diffStage_controlPipe_payload_lastRow) begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_144[7:0];
                    end else begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_146[7:0];
                    end
                  end else begin
                    if(diffStage_controlPipe_payload_lastRow) begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_148[7:0];
                    end else begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_150[7:0];
                    end
                  end
                end else begin
                  if(when_SuperResolutionPart3_l1009) begin
                    if(diffStage_controlPipe_payload_lastRow) begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_152[7:0];
                    end else begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_154[7:0];
                    end
                  end else begin
                    if(diffStage_controlPipe_payload_lastRow) begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_156[7:0];
                    end else begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_158[7:0];
                    end
                  end
                end
              end
            end
          end else begin
            if(when_SuperResolutionPart3_l1018) begin
              if(when_SuperResolutionPart3_l1019) begin
                if(when_SuperResolutionPart3_l1020) begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_160[7:0];
                end else begin
                  if(when_SuperResolutionPart3_l1021) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_162[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_164[7:0];
                  end
                end
              end else begin
                if(when_SuperResolutionPart3_l1024) begin
                  if(when_SuperResolutionPart3_l1025) begin
                    if(diffStage_controlPipe_payload_firstRow) begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_166[7:0];
                    end else begin
                      if(diffStage_controlPipe_payload_lastRow) begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_168[7:0];
                      end else begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_170[7:0];
                      end
                    end
                  end else begin
                    if(diffStage_controlPipe_payload_lastRow) begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_172[7:0];
                    end else begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_174[7:0];
                    end
                  end
                end else begin
                  if(when_SuperResolutionPart3_l1033) begin
                    if(when_SuperResolutionPart3_l1034) begin
                      if(diffStage_controlPipe_payload_lastRow) begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_176[7:0];
                      end else begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_178[7:0];
                      end
                    end else begin
                      if(diffStage_controlPipe_payload_lastRow) begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_180[7:0];
                      end else begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_182[7:0];
                      end
                    end
                  end else begin
                    if(when_SuperResolutionPart3_l1042) begin
                      if(diffStage_controlPipe_payload_lastRow) begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_184[7:0];
                      end else begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_186[7:0];
                      end
                    end else begin
                      if(diffStage_controlPipe_payload_lastRow) begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_188[7:0];
                      end else begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_190[7:0];
                      end
                    end
                  end
                end
              end
            end else begin
              if(when_SuperResolutionPart3_l1051) begin
                if(when_SuperResolutionPart3_l1052) begin
                  if(when_SuperResolutionPart3_l1053) begin
                    if(diffStage_controlPipe_payload_firstRow) begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_192[7:0];
                    end else begin
                      if(diffStage_controlPipe_payload_lastRow) begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_194[7:0];
                      end else begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_196[7:0];
                      end
                    end
                  end else begin
                    if(diffStage_controlPipe_payload_lastRow) begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_198[7:0];
                    end else begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_200[7:0];
                    end
                  end
                end else begin
                  if(when_SuperResolutionPart3_l1061) begin
                    if(when_SuperResolutionPart3_l1062) begin
                      if(diffStage_controlPipe_payload_lastRow) begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_202[7:0];
                      end else begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_204[7:0];
                      end
                    end else begin
                      if(diffStage_controlPipe_payload_lastRow) begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_206[7:0];
                      end else begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_208[7:0];
                      end
                    end
                  end else begin
                    if(when_SuperResolutionPart3_l1070) begin
                      if(diffStage_controlPipe_payload_lastRow) begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_210[7:0];
                      end else begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_212[7:0];
                      end
                    end else begin
                      if(diffStage_controlPipe_payload_lastRow) begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_214[7:0];
                      end else begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_216[7:0];
                      end
                    end
                  end
                end
              end else begin
                if(when_SuperResolutionPart3_l1078) begin
                  if(when_SuperResolutionPart3_l1079) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_218[7:0];
                  end else begin
                    if(when_SuperResolutionPart3_l1080) begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_220[7:0];
                    end else begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_222[7:0];
                    end
                  end
                end else begin
                  if(when_SuperResolutionPart3_l1082) begin
                    if(when_SuperResolutionPart3_l1083) begin
                      if(when_SuperResolutionPart3_l1084) begin
                        if(diffStage_controlPipe_payload_firstRow) begin
                          resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_224[7:0];
                        end else begin
                          if(diffStage_controlPipe_payload_lastRow) begin
                            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_226[7:0];
                          end else begin
                            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_228[7:0];
                          end
                        end
                      end else begin
                        if(diffStage_controlPipe_payload_lastRow) begin
                          resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_230[7:0];
                        end else begin
                          resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_232[7:0];
                        end
                      end
                    end else begin
                      if(when_SuperResolutionPart3_l1092) begin
                        if(when_SuperResolutionPart3_l1093) begin
                          if(diffStage_controlPipe_payload_lastRow) begin
                            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_234[7:0];
                          end else begin
                            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_236[7:0];
                          end
                        end else begin
                          if(diffStage_controlPipe_payload_lastRow) begin
                            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_238[7:0];
                          end else begin
                            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_240[7:0];
                          end
                        end
                      end else begin
                        if(when_SuperResolutionPart3_l1101) begin
                          if(diffStage_controlPipe_payload_lastRow) begin
                            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_242[7:0];
                          end else begin
                            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_244[7:0];
                          end
                        end else begin
                          if(diffStage_controlPipe_payload_lastRow) begin
                            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_246[7:0];
                          end else begin
                            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_248[7:0];
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
  end

  assign when_SuperResolutionPart3_l840 = ((diffStage_controlPipe_payload_currentPosition == 2'b00) && diffStage_mainOneValidStream_payload);
  assign when_SuperResolutionPart3_l846 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l847 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l850 = (minDiff < diffStage_controlPipe_payload_verticalDiff);
  assign when_SuperResolutionPart3_l854 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l855 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l860 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l861 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l851 = (diffStage_controlPipe_payload_verticalDiff == minDiff);
  assign when_SuperResolutionPart3_l841 = ((diffStage_controlPipe_payload_currentPosition == 2'b01) && diffStage_mainTwoValidStream_payload);
  assign when_SuperResolutionPart3_l842 = ((diffStage_controlPipe_payload_currentPosition == 2'b10) && diffStage_mainThreeValidStream_payload);
  assign when_SuperResolutionPart3_l869 = ((diffStage_controlPipe_payload_horizontalDirectionValid && diffStage_controlPipe_payload_mainDirectionValid) && diffStage_controlPipe_payload_counterDirectionValid);
  assign when_SuperResolutionPart3_l870 = ((diffStage_controlPipe_payload_horizontalDiff <= diffStage_controlPipe_payload_mainDiff) && (diffStage_controlPipe_payload_horizontalDiff <= diffStage_controlPipe_payload_counterDiff));
  assign when_SuperResolutionPart3_l871 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l872 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l875 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l876 = (diffStage_controlPipe_payload_nextPosition == 2'b01);
  assign when_SuperResolutionPart3_l885 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l893 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l884 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l902 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l903 = (diffStage_controlPipe_payload_nextPosition == 2'b01);
  assign when_SuperResolutionPart3_l912 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l920 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l911 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l874 = ((diffStage_controlPipe_payload_mainDiff < diffStage_controlPipe_payload_horizontalDiff) && (diffStage_controlPipe_payload_mainDiff <= diffStage_controlPipe_payload_counterDiff));
  assign when_SuperResolutionPart3_l930 = (diffStage_controlPipe_payload_mainDiff <= diffStage_controlPipe_payload_counterDiff);
  assign when_SuperResolutionPart3_l931 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l932 = (diffStage_controlPipe_payload_nextPosition == 2'b01);
  assign when_SuperResolutionPart3_l941 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l949 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l940 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l958 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l959 = (diffStage_controlPipe_payload_nextPosition == 2'b01);
  assign when_SuperResolutionPart3_l968 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l976 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l967 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l986 = (diffStage_controlPipe_payload_horizontalDiff <= diffStage_controlPipe_payload_counterDiff);
  assign when_SuperResolutionPart3_l987 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l988 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l991 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l992 = (diffStage_controlPipe_payload_nextPosition == 2'b01);
  assign when_SuperResolutionPart3_l1001 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l1009 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l1000 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l1019 = (diffStage_controlPipe_payload_horizontalDiff <= diffStage_controlPipe_payload_mainDiff);
  assign when_SuperResolutionPart3_l1020 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l1021 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l1024 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l1025 = (diffStage_controlPipe_payload_nextPosition == 2'b01);
  assign when_SuperResolutionPart3_l1034 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l1042 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l1033 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l1052 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l1053 = (diffStage_controlPipe_payload_nextPosition == 2'b01);
  assign when_SuperResolutionPart3_l1062 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l1070 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l1061 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l1079 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l1080 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l1083 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l1084 = (diffStage_controlPipe_payload_nextPosition == 2'b01);
  assign when_SuperResolutionPart3_l1093 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l1101 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l1092 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l929 = (((! diffStage_controlPipe_payload_horizontalDirectionValid) && diffStage_controlPipe_payload_mainDirectionValid) && diffStage_controlPipe_payload_counterDirectionValid);
  assign when_SuperResolutionPart3_l985 = ((diffStage_controlPipe_payload_horizontalDirectionValid && (! diffStage_controlPipe_payload_mainDirectionValid)) && diffStage_controlPipe_payload_counterDirectionValid);
  assign when_SuperResolutionPart3_l1018 = ((diffStage_controlPipe_payload_horizontalDirectionValid && diffStage_controlPipe_payload_mainDirectionValid) && (! diffStage_controlPipe_payload_counterDirectionValid));
  assign when_SuperResolutionPart3_l1051 = (((! diffStage_controlPipe_payload_horizontalDirectionValid) && (! diffStage_controlPipe_payload_mainDirectionValid)) && diffStage_controlPipe_payload_counterDirectionValid);
  assign when_SuperResolutionPart3_l1078 = ((diffStage_controlPipe_payload_horizontalDirectionValid && (! diffStage_controlPipe_payload_mainDirectionValid)) && (! diffStage_controlPipe_payload_counterDirectionValid));
  assign when_SuperResolutionPart3_l1082 = (((! diffStage_controlPipe_payload_horizontalDirectionValid) && diffStage_controlPipe_payload_mainDirectionValid) && (! diffStage_controlPipe_payload_counterDirectionValid));
  assign resultStage_pixelStream_ready = (! resultStage_pixelStream_rValid);
  assign resultStage_pixelStream_s2mPipe_valid = (resultStage_pixelStream_valid || resultStage_pixelStream_rValid);
  assign resultStage_pixelStream_s2mPipe_payload = (resultStage_pixelStream_rValid ? resultStage_pixelStream_rData : resultStage_pixelStream_payload);
  always @(*) begin
    resultStage_pixelStream_s2mPipe_ready = resultStage_resultStream_ready;
    if(when_Stream_l368_67) begin
      resultStage_pixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_67 = (! resultStage_resultStream_valid);
  assign resultStage_resultStream_valid = resultStage_pixelStream_s2mPipe_rValid;
  assign resultStage_resultStream_payload = resultStage_pixelStream_s2mPipe_rData;
  assign when_SuperResolutionPart3_l1115 = (! resultStage_controlPipeBeforePipe_payload_finalResult);
  assign diffStage_controlPipe_fire = (diffStage_controlPipe_valid && diffStage_controlPipe_ready);
  assign CICC1851_resultStage_mainOnePixelStream_ready_2 = (CICC1851_resultStage_mainOnePixelStream_ready && CICC1851_resultStage_mainOnePixelStream_ready_1);
  assign CICC1851_resultStage_mainOnePixelStream_ready = (((((((((((((resultStage_resultStream_valid && resultStage_mainOnePixelStream_valid) && resultStage_counterOnePixelStream_valid) && resultStage_mainTwoPixelStream_valid) && resultStage_counterTwoPixelStream_valid) && resultStage_mainThreePixelStream_valid) && resultStage_counterThreePixelStream_valid) && resultStage_mainOneValidStream_valid) && resultStage_counterOneValidStream_valid) && resultStage_mainTwoValidStream_valid) && resultStage_counterTwoValidStream_valid) && resultStage_mainThreeValidStream_valid) && resultStage_counterThreeValidStream_valid) && resultStage_controlPipe_valid);
  assign resultStage_resultStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_mainOnePixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_counterOnePixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_mainTwoPixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_counterTwoPixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_mainThreePixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_counterThreePixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_mainOneValidStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_counterOneValidStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_mainTwoValidStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_counterTwoValidStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_mainThreeValidStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_counterThreeValidStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_controlPipe_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign when_Stream_l438 = ((! resultStage_controlPipe_payload_pipeValid) || (! resultStage_controlPipe_payload_finalResult));
  always @(*) begin
    resultsJoin_valid = CICC1851_resultStage_mainOnePixelStream_ready;
    if(when_Stream_l438) begin
      resultsJoin_valid = 1'b0;
    end
  end

  always @(*) begin
    CICC1851_resultStage_mainOnePixelStream_ready_1 = resultsJoin_ready;
    if(when_Stream_l438) begin
      CICC1851_resultStage_mainOnePixelStream_ready_1 = 1'b1;
    end
  end

  assign pixelsStream_valid = resultsJoin_valid;
  assign resultsJoin_ready = pixelsStream_ready;
  assign pixelsStream_payload_pixel = resultStage_resultStream_payload;
  assign pixelsStream_payload_frameStart = resultStage_controlPipe_payload_frameStart;
  assign pixelsStream_payload_rowEnd = resultStage_controlPipe_payload_rowEnd;
  assign pixelsStream_ready = (! pixelsStream_rValid);
  assign pixelsStream_s2mPipe_valid = (pixelsStream_valid || pixelsStream_rValid);
  assign pixelsStream_s2mPipe_payload_pixel = (pixelsStream_rValid ? pixelsStream_rData_pixel : pixelsStream_payload_pixel);
  assign pixelsStream_s2mPipe_payload_frameStart = (pixelsStream_rValid ? pixelsStream_rData_frameStart : pixelsStream_payload_frameStart);
  assign pixelsStream_s2mPipe_payload_rowEnd = (pixelsStream_rValid ? pixelsStream_rData_rowEnd : pixelsStream_payload_rowEnd);
  always @(*) begin
    pixelsStream_s2mPipe_ready = pixelsStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_68) begin
      pixelsStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_68 = (! pixelsStream_s2mPipe_m2sPipe_valid);
  assign pixelsStream_s2mPipe_m2sPipe_valid = pixelsStream_s2mPipe_rValid;
  assign pixelsStream_s2mPipe_m2sPipe_payload_pixel = pixelsStream_s2mPipe_rData_pixel;
  assign pixelsStream_s2mPipe_m2sPipe_payload_frameStart = pixelsStream_s2mPipe_rData_frameStart;
  assign pixelsStream_s2mPipe_m2sPipe_payload_rowEnd = pixelsStream_s2mPipe_rData_rowEnd;
  assign pixelsStream_s2mPipe_m2sPipe_ready = pixelsOut_ready;
  assign controlStateMachine_wantExit = 1'b0;
  always @(*) begin
    controlStateMachine_wantStart = 1'b0;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_8_HOLD : begin
      end
      controlStateMachine_enumDef_8_PASS : begin
      end
      controlStateMachine_enumDef_8_EXTRA : begin
      end
      default : begin
        controlStateMachine_wantStart = 1'b1;
      end
    endcase
  end

  assign controlStateMachine_wantKill = 1'b0;
  always @(*) begin
    controlStateMachine_stateNext = controlStateMachine_stateReg;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_8_HOLD : begin
        if(passPixels_fire_13) begin
          if(when_SuperResolutionPart3_l1158) begin
            controlStateMachine_stateNext = controlStateMachine_enumDef_8_PASS;
          end
        end
      end
      controlStateMachine_enumDef_8_PASS : begin
        if(controlStream_fire) begin
          controlStateMachine_stateNext = controlStateMachine_enumDef_8_EXTRA;
        end
      end
      controlStateMachine_enumDef_8_EXTRA : begin
        if(controlStream_fire_1) begin
          if(writeDone) begin
            if(when_SuperResolutionPart3_l1199) begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_8_HOLD;
            end else begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_8_PASS;
            end
          end else begin
            if(outReachRowEnd) begin
              if(when_SuperResolutionPart3_l1202) begin
                controlStateMachine_stateNext = controlStateMachine_enumDef_8_PASS;
              end else begin
                controlStateMachine_stateNext = controlStateMachine_enumDef_8_HOLD;
              end
            end else begin
              if(when_SuperResolutionPart3_l1205) begin
                controlStateMachine_stateNext = controlStateMachine_enumDef_8_PASS;
              end else begin
                controlStateMachine_stateNext = controlStateMachine_enumDef_8_HOLD;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
    if(controlStateMachine_wantStart) begin
      controlStateMachine_stateNext = controlStateMachine_enumDef_8_HOLD;
    end
    if(controlStateMachine_wantKill) begin
      controlStateMachine_stateNext = controlStateMachine_enumDef_8_BOOT;
    end
  end

  assign passPixels_fire_13 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart3_l1158 = ((outRowCount_value < bufferRowCount_value) && (outPixelAddr_value < bufferWAddr_value));
  assign controlStream_fire = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart3_l1168 = (outPixelAddr_value == 12'h0);
  assign when_SuperResolutionPart3_l1188 = (outRowCount_value == 12'h0);
  assign controlStream_fire_1 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart3_l1199 = (outReachFinalRow && outReachRowEnd);
  assign passPixels_fire_14 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart3_l1202 = (((bufferRowCount_value == CICC1851_when_SuperResolutionPart3_l1202) || (12'h001 < bufferWAddr_value)) || ((bufferWAddr_value == 12'h001) && passPixels_fire_14));
  assign passPixels_fire_15 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart3_l1205 = (((CICC1851_when_SuperResolutionPart3_l1205 < bufferRowCount_value) || ((bufferWAddr_value == CICC1851_when_SuperResolutionPart3_l1205_1) && passPixels_fire_15)) || (CICC1851_when_SuperResolutionPart3_l1205_2 < bufferWAddr_value));
  assign when_SuperResolutionPart3_l1217 = (outRowCount_value == 12'h0);
  assign controlStream_fire_2 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart3_l1220 = (frameStart && controlStream_fire_2);
  assign controlStream_fire_3 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart3_l1223 = (controlStream_fire_3 && (CICC1851_when_SuperResolutionPart3_l1223 == CICC1851_when_SuperResolutionPart3_l1223_1));
  assign controlStream_fire_4 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart3_l1224 = ((outReachRowEnd && (CICC1851_when_SuperResolutionPart3_l1224 == CICC1851_when_SuperResolutionPart3_l1224_1)) && controlStream_fire_4);
  assign controlStream_fire_5 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart3_l1226 = (controlStream_fire_5 && outReachRowEnd);
  assign controlStream_fire_6 = (controlStream_valid && controlStream_ready);
  assign controlStream_fire_7 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart3_l1247 = (controlStream_payload_rowEnd && controlStream_fire_7);
  assign when_SuperResolutionPart3_l1248 = (outRowCount_value != 12'h0);
  assign when_SuperResolutionPart3_l1250 = (currentRowBuffer == 2'b10);
  assign when_SuperResolutionPart3_l1252 = (nextRowBuffer == 2'b10);
  always @(posedge clk or negedge resetn) begin
    if(!resetn) begin
      inpThreeDone <= 1'b0;
      readDone <= 1'b0;
      startRead <= 1'b0;
      frameStart <= 1'b0;
      inpThreshold <= 8'h80;
      bmpWidth <= 10'h3c0;
      bmpHeight <= 10'h21c;
      holdBuffer <= 1'b0;
      writeDone <= 1'b0;
      bufferRowCount_value <= 12'h0;
      bufferEnable <= 1'b0;
      bufferSwitch <= 2'b00;
      nextRowBuffer <= 2'b01;
      currentRowBuffer <= 2'b00;
      bufferReuse <= 1'b0;
      bufferWAddr_value <= 12'h0;
      outPixelAddr_value <= 12'h0;
      outRowCount_value <= 12'h0;
      alreadySendRow_value <= 12'h0;
      alreadySendCountInRow_value <= 12'h0;
      alreadyReachRowEnd <= 1'b0;
      alreadyReachFinalRow <= 1'b0;
      outReachRowEnd <= 1'b0;
      outReachFinalRow <= 1'b0;
      bufferReachRowEnd <= 1'b0;
      bufferReachFinalRow <= 1'b0;
      minDiff <= 8'h0;
      candidatePixel <= 8'h0;
      isHorizontalDirection <= 1'b0;
      inValidMinDiff <= 1'b0;
      pixelsIn_rValid <= 1'b0;
      pixelsIn_s2mPipe_rValid <= 1'b0;
      mainPixelAddrOneStream_rValid <= 1'b0;
      mainPixelAddrOneStream_s2mPipe_rValid <= 1'b0;
      CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_mainOnePixelStream_valid <= 1'b0;
      counterPixelAddrOneStream_rValid <= 1'b0;
      counterPixelAddrOneStream_s2mPipe_rValid <= 1'b0;
      CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_counterOnePixelStream_valid <= 1'b0;
      mainPixelAddrTwoStream_rValid <= 1'b0;
      mainPixelAddrTwoStream_s2mPipe_rValid <= 1'b0;
      CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_mainTwoPixelStream_valid <= 1'b0;
      counterPixelAddrTwoStream_rValid <= 1'b0;
      counterPixelAddrTwoStream_s2mPipe_rValid <= 1'b0;
      CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_counterTwoPixelStream_valid <= 1'b0;
      mainPixelAddrThreeStream_rValid <= 1'b0;
      mainPixelAddrThreeStream_s2mPipe_rValid <= 1'b0;
      CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_mainThreePixelStream_valid <= 1'b0;
      counterPixelAddrThreeStream_rValid <= 1'b0;
      counterPixelAddrThreeStream_s2mPipe_rValid <= 1'b0;
      CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_counterThreePixelStream_valid <= 1'b0;
      mainValidAddrOneStream_rValid <= 1'b0;
      mainValidAddrOneStream_s2mPipe_rValid <= 1'b0;
      CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_mainOneValidStream_valid <= 1'b0;
      counterValidAddrOneStream_rValid <= 1'b0;
      counterValidAddrOneStream_s2mPipe_rValid <= 1'b0;
      CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_counterOneValidStream_valid <= 1'b0;
      mainValidAddrTwoStream_rValid <= 1'b0;
      mainValidAddrTwoStream_s2mPipe_rValid <= 1'b0;
      CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_mainTwoValidStream_valid <= 1'b0;
      counterValidAddrTwoStream_rValid <= 1'b0;
      counterValidAddrTwoStream_s2mPipe_rValid <= 1'b0;
      CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_counterTwoValidStream_valid <= 1'b0;
      mainValidAddrThreeStream_rValid <= 1'b0;
      mainValidAddrThreeStream_s2mPipe_rValid <= 1'b0;
      CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_mainThreeValidStream_valid <= 1'b0;
      counterValidAddrThreeStream_rValid <= 1'b0;
      counterValidAddrThreeStream_s2mPipe_rValid <= 1'b0;
      CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_counterThreeValidStream_valid <= 1'b0;
      controlStream_rValid <= 1'b0;
      controlStream_s2mPipe_rValid <= 1'b0;
      controlStream_s2mPipe_m2sPipe_rValid <= 1'b0;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rValid <= 1'b0;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rValid <= 1'b0;
      readStage_mainOnePixelStream_rValid <= 1'b0;
      readStage_mainOnePixelStream_s2mPipe_rValid <= 1'b0;
      readStage_counterOnePixelStream_rValid <= 1'b0;
      readStage_counterOnePixelStream_s2mPipe_rValid <= 1'b0;
      readStage_mainTwoPixelStream_rValid <= 1'b0;
      readStage_mainTwoPixelStream_s2mPipe_rValid <= 1'b0;
      readStage_counterTwoPixelStream_rValid <= 1'b0;
      readStage_counterTwoPixelStream_s2mPipe_rValid <= 1'b0;
      readStage_mainThreePixelStream_rValid <= 1'b0;
      readStage_mainThreePixelStream_s2mPipe_rValid <= 1'b0;
      readStage_counterThreePixelStream_rValid <= 1'b0;
      readStage_counterThreePixelStream_s2mPipe_rValid <= 1'b0;
      readStage_mainOneValidStream_rValid <= 1'b0;
      readStage_mainOneValidStream_s2mPipe_rValid <= 1'b0;
      readStage_counterOneValidStream_rValid <= 1'b0;
      readStage_counterOneValidStream_s2mPipe_rValid <= 1'b0;
      readStage_mainTwoValidStream_rValid <= 1'b0;
      readStage_mainTwoValidStream_s2mPipe_rValid <= 1'b0;
      readStage_counterTwoValidStream_rValid <= 1'b0;
      readStage_counterTwoValidStream_s2mPipe_rValid <= 1'b0;
      readStage_mainThreeValidStream_rValid <= 1'b0;
      readStage_mainThreeValidStream_s2mPipe_rValid <= 1'b0;
      readStage_counterThreeValidStream_rValid <= 1'b0;
      readStage_counterThreeValidStream_s2mPipe_rValid <= 1'b0;
      readStage_controlPipe_translated_rValid <= 1'b0;
      readStage_controlPipe_translated_s2mPipe_rValid <= 1'b0;
      compareStage_mainOnePixelStream_rValid <= 1'b0;
      compareStage_mainOnePixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_counterOnePixelStream_rValid <= 1'b0;
      compareStage_counterOnePixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_mainTwoPixelStream_rValid <= 1'b0;
      compareStage_mainTwoPixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_counterTwoPixelStream_rValid <= 1'b0;
      compareStage_counterTwoPixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_mainThreePixelStream_rValid <= 1'b0;
      compareStage_mainThreePixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_counterThreePixelStream_rValid <= 1'b0;
      compareStage_counterThreePixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_mainOneValidStream_rValid <= 1'b0;
      compareStage_mainOneValidStream_s2mPipe_rValid <= 1'b0;
      compareStage_counterOneValidStream_rValid <= 1'b0;
      compareStage_counterOneValidStream_s2mPipe_rValid <= 1'b0;
      compareStage_mainTwoValidStream_rValid <= 1'b0;
      compareStage_mainTwoValidStream_s2mPipe_rValid <= 1'b0;
      compareStage_counterTwoValidStream_rValid <= 1'b0;
      compareStage_counterTwoValidStream_s2mPipe_rValid <= 1'b0;
      compareStage_mainThreeValidStream_rValid <= 1'b0;
      compareStage_mainThreeValidStream_s2mPipe_rValid <= 1'b0;
      compareStage_counterThreeValidStream_rValid <= 1'b0;
      compareStage_counterThreeValidStream_s2mPipe_rValid <= 1'b0;
      compareStage_controlPipe_translated_rValid <= 1'b0;
      compareStage_controlPipe_translated_s2mPipe_rValid <= 1'b0;
      diffStage_mainOnePixelStream_rValid <= 1'b0;
      diffStage_mainOnePixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_counterOnePixelStream_rValid <= 1'b0;
      diffStage_counterOnePixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_mainTwoPixelStream_rValid <= 1'b0;
      diffStage_mainTwoPixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_counterTwoPixelStream_rValid <= 1'b0;
      diffStage_counterTwoPixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_mainThreePixelStream_rValid <= 1'b0;
      diffStage_mainThreePixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_counterThreePixelStream_rValid <= 1'b0;
      diffStage_counterThreePixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_mainOneValidStream_rValid <= 1'b0;
      diffStage_mainOneValidStream_s2mPipe_rValid <= 1'b0;
      diffStage_counterOneValidStream_rValid <= 1'b0;
      diffStage_counterOneValidStream_s2mPipe_rValid <= 1'b0;
      diffStage_mainTwoValidStream_rValid <= 1'b0;
      diffStage_mainTwoValidStream_s2mPipe_rValid <= 1'b0;
      diffStage_counterTwoValidStream_rValid <= 1'b0;
      diffStage_counterTwoValidStream_s2mPipe_rValid <= 1'b0;
      diffStage_mainThreeValidStream_rValid <= 1'b0;
      diffStage_mainThreeValidStream_s2mPipe_rValid <= 1'b0;
      diffStage_counterThreeValidStream_rValid <= 1'b0;
      diffStage_counterThreeValidStream_s2mPipe_rValid <= 1'b0;
      resultStage_controlPipeBeforePipe_rValid <= 1'b0;
      resultStage_controlPipeBeforePipe_s2mPipe_rValid <= 1'b0;
      resultStage_pixelStream_rValid <= 1'b0;
      resultStage_pixelStream_s2mPipe_rValid <= 1'b0;
      pixelsStream_rValid <= 1'b0;
      pixelsStream_s2mPipe_rValid <= 1'b0;
      controlStateMachine_stateReg <= controlStateMachine_enumDef_8_BOOT;
    end else begin
      if(when_SuperResolutionPart3_l72) begin
        inpThreeDone <= 1'b0;
      end
      if(when_SuperResolutionPart3_l75) begin
        readDone <= 1'b0;
      end
      if(when_SuperResolutionPart3_l78) begin
        startRead <= 1'b1;
      end
      if(when_SuperResolutionPart3_l78_1) begin
        startRead <= 1'b0;
      end
      inpThreshold <= thresholdIn;
      bmpWidth <= widthIn;
      bmpHeight <= heightIn;
      if(when_SuperResolutionPart3_l93) begin
        holdBuffer <= 1'b0;
      end
      if(when_SuperResolutionPart3_l96) begin
        writeDone <= 1'b0;
      end
      bufferRowCount_value <= bufferRowCount_valueNext;
      if(when_SuperResolutionPart3_l102) begin
        bufferEnable <= 1'b1;
      end
      if(when_SuperResolutionPart3_l102_1) begin
        bufferEnable <= 1'b0;
      end
      if(inpThreeDone) begin
        bufferReuse <= 1'b0;
      end
      bufferWAddr_value <= bufferWAddr_valueNext;
      outPixelAddr_value <= outPixelAddr_valueNext;
      outRowCount_value <= outRowCount_valueNext;
      alreadySendRow_value <= alreadySendRow_valueNext;
      alreadySendCountInRow_value <= alreadySendCountInRow_valueNext;
      if(when_SuperResolutionPart3_l154) begin
        bufferSwitch <= 2'b00;
        nextRowBuffer <= {1'd0, CICC1851_nextRowBuffer};
        currentRowBuffer <= 2'b00;
        minDiff <= 8'h0;
        candidatePixel <= 8'h0;
        isHorizontalDirection <= 1'b0;
      end
      if(pixelsIn_valid) begin
        pixelsIn_rValid <= 1'b1;
      end
      if(pixelsIn_s2mPipe_ready) begin
        pixelsIn_rValid <= 1'b0;
      end
      if(pixelsIn_s2mPipe_ready) begin
        pixelsIn_s2mPipe_rValid <= pixelsIn_s2mPipe_valid;
      end
      if(when_SuperResolutionPart3_l226) begin
        bufferReachRowEnd <= 1'b1;
      end
      if(when_SuperResolutionPart3_l227) begin
        bufferReachFinalRow <= 1'b1;
      end
      if(when_SuperResolutionPart3_l230) begin
        if(bufferReachFinalRow) begin
          bufferReuse <= 1'b1;
          bufferReachRowEnd <= 1'b0;
          bufferReachFinalRow <= 1'b0;
        end else begin
          bufferReachRowEnd <= 1'b0;
        end
      end
      if(when_SuperResolutionPart3_l243) begin
        if(when_SuperResolutionPart3_l244) begin
          bufferSwitch <= 2'b00;
        end else begin
          bufferSwitch <= (bufferSwitch + 2'b01);
        end
      end
      if(when_SuperResolutionPart3_l251) begin
        holdBuffer <= 1'b1;
        bufferEnable <= 1'b0;
        if(when_SuperResolutionPart3_l255) begin
          writeDone <= 1'b1;
          bufferEnable <= 1'b0;
        end
      end
      if(when_SuperResolutionPart3_l262) begin
        frameStart <= 1'b1;
      end
      if(inpThreeDone) begin
        inpThreeDone <= 1'b0;
      end
      if(when_SuperResolutionPart3_l270) begin
        alreadyReachRowEnd <= 1'b1;
      end
      if(when_SuperResolutionPart3_l271) begin
        alreadyReachFinalRow <= 1'b1;
      end
      if(pixelsOut_fire_2) begin
        if(alreadyReachRowEnd) begin
          alreadyReachRowEnd <= 1'b0;
          if(alreadyReachFinalRow) begin
            alreadyReachFinalRow <= 1'b0;
          end
        end
      end
      if(when_SuperResolutionPart3_l282) begin
        inpThreeDone <= 1'b1;
      end
      if(mainPixelAddrOneStream_valid) begin
        mainPixelAddrOneStream_rValid <= 1'b1;
      end
      if(mainPixelAddrOneStream_s2mPipe_ready) begin
        mainPixelAddrOneStream_rValid <= 1'b0;
      end
      if(mainPixelAddrOneStream_s2mPipe_ready) begin
        mainPixelAddrOneStream_s2mPipe_rValid <= mainPixelAddrOneStream_s2mPipe_valid;
      end
      if(CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(mainPixelAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_2 <= mainPixelAddrOneStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_1) begin
        CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_1) begin
        CICC1851_readStage_mainOnePixelStream_valid <= (CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready || CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_3);
      end
      if(counterPixelAddrOneStream_valid) begin
        counterPixelAddrOneStream_rValid <= 1'b1;
      end
      if(counterPixelAddrOneStream_s2mPipe_ready) begin
        counterPixelAddrOneStream_rValid <= 1'b0;
      end
      if(counterPixelAddrOneStream_s2mPipe_ready) begin
        counterPixelAddrOneStream_s2mPipe_rValid <= counterPixelAddrOneStream_s2mPipe_valid;
      end
      if(CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(counterPixelAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_2 <= counterPixelAddrOneStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_2) begin
        CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_2) begin
        CICC1851_readStage_counterOnePixelStream_valid <= (CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready || CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_3);
      end
      if(mainPixelAddrTwoStream_valid) begin
        mainPixelAddrTwoStream_rValid <= 1'b1;
      end
      if(mainPixelAddrTwoStream_s2mPipe_ready) begin
        mainPixelAddrTwoStream_rValid <= 1'b0;
      end
      if(mainPixelAddrTwoStream_s2mPipe_ready) begin
        mainPixelAddrTwoStream_s2mPipe_rValid <= mainPixelAddrTwoStream_s2mPipe_valid;
      end
      if(CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= mainPixelAddrTwoStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_3) begin
        CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_3) begin
        CICC1851_readStage_mainTwoPixelStream_valid <= (CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready || CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_3);
      end
      if(counterPixelAddrTwoStream_valid) begin
        counterPixelAddrTwoStream_rValid <= 1'b1;
      end
      if(counterPixelAddrTwoStream_s2mPipe_ready) begin
        counterPixelAddrTwoStream_rValid <= 1'b0;
      end
      if(counterPixelAddrTwoStream_s2mPipe_ready) begin
        counterPixelAddrTwoStream_s2mPipe_rValid <= counterPixelAddrTwoStream_s2mPipe_valid;
      end
      if(CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= counterPixelAddrTwoStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_4) begin
        CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_4) begin
        CICC1851_readStage_counterTwoPixelStream_valid <= (CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready || CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_3);
      end
      if(mainPixelAddrThreeStream_valid) begin
        mainPixelAddrThreeStream_rValid <= 1'b1;
      end
      if(mainPixelAddrThreeStream_s2mPipe_ready) begin
        mainPixelAddrThreeStream_rValid <= 1'b0;
      end
      if(mainPixelAddrThreeStream_s2mPipe_ready) begin
        mainPixelAddrThreeStream_s2mPipe_rValid <= mainPixelAddrThreeStream_s2mPipe_valid;
      end
      if(CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_2 <= mainPixelAddrThreeStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_5) begin
        CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_5) begin
        CICC1851_readStage_mainThreePixelStream_valid <= (CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready || CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_3);
      end
      if(counterPixelAddrThreeStream_valid) begin
        counterPixelAddrThreeStream_rValid <= 1'b1;
      end
      if(counterPixelAddrThreeStream_s2mPipe_ready) begin
        counterPixelAddrThreeStream_rValid <= 1'b0;
      end
      if(counterPixelAddrThreeStream_s2mPipe_ready) begin
        counterPixelAddrThreeStream_s2mPipe_rValid <= counterPixelAddrThreeStream_s2mPipe_valid;
      end
      if(CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_2 <= counterPixelAddrThreeStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_6) begin
        CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_6) begin
        CICC1851_readStage_counterThreePixelStream_valid <= (CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready || CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_3);
      end
      if(mainValidAddrOneStream_valid) begin
        mainValidAddrOneStream_rValid <= 1'b1;
      end
      if(mainValidAddrOneStream_s2mPipe_ready) begin
        mainValidAddrOneStream_rValid <= 1'b0;
      end
      if(mainValidAddrOneStream_s2mPipe_ready) begin
        mainValidAddrOneStream_s2mPipe_rValid <= mainValidAddrOneStream_s2mPipe_valid;
      end
      if(CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(mainValidAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_2 <= mainValidAddrOneStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_7) begin
        CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_7) begin
        CICC1851_readStage_mainOneValidStream_valid <= (CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready || CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_3);
      end
      if(counterValidAddrOneStream_valid) begin
        counterValidAddrOneStream_rValid <= 1'b1;
      end
      if(counterValidAddrOneStream_s2mPipe_ready) begin
        counterValidAddrOneStream_rValid <= 1'b0;
      end
      if(counterValidAddrOneStream_s2mPipe_ready) begin
        counterValidAddrOneStream_s2mPipe_rValid <= counterValidAddrOneStream_s2mPipe_valid;
      end
      if(CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(counterValidAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_2 <= counterValidAddrOneStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_8) begin
        CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_8) begin
        CICC1851_readStage_counterOneValidStream_valid <= (CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready || CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_3);
      end
      if(mainValidAddrTwoStream_valid) begin
        mainValidAddrTwoStream_rValid <= 1'b1;
      end
      if(mainValidAddrTwoStream_s2mPipe_ready) begin
        mainValidAddrTwoStream_rValid <= 1'b0;
      end
      if(mainValidAddrTwoStream_s2mPipe_ready) begin
        mainValidAddrTwoStream_s2mPipe_rValid <= mainValidAddrTwoStream_s2mPipe_valid;
      end
      if(CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(mainValidAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= mainValidAddrTwoStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_9) begin
        CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_9) begin
        CICC1851_readStage_mainTwoValidStream_valid <= (CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready || CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_3);
      end
      if(counterValidAddrTwoStream_valid) begin
        counterValidAddrTwoStream_rValid <= 1'b1;
      end
      if(counterValidAddrTwoStream_s2mPipe_ready) begin
        counterValidAddrTwoStream_rValid <= 1'b0;
      end
      if(counterValidAddrTwoStream_s2mPipe_ready) begin
        counterValidAddrTwoStream_s2mPipe_rValid <= counterValidAddrTwoStream_s2mPipe_valid;
      end
      if(CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(counterValidAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= counterValidAddrTwoStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_10) begin
        CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_10) begin
        CICC1851_readStage_counterTwoValidStream_valid <= (CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready || CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_3);
      end
      if(mainValidAddrThreeStream_valid) begin
        mainValidAddrThreeStream_rValid <= 1'b1;
      end
      if(mainValidAddrThreeStream_s2mPipe_ready) begin
        mainValidAddrThreeStream_rValid <= 1'b0;
      end
      if(mainValidAddrThreeStream_s2mPipe_ready) begin
        mainValidAddrThreeStream_s2mPipe_rValid <= mainValidAddrThreeStream_s2mPipe_valid;
      end
      if(CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(mainValidAddrThreeStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_2 <= mainValidAddrThreeStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_11) begin
        CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_11) begin
        CICC1851_readStage_mainThreeValidStream_valid <= (CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready || CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_3);
      end
      if(counterValidAddrThreeStream_valid) begin
        counterValidAddrThreeStream_rValid <= 1'b1;
      end
      if(counterValidAddrThreeStream_s2mPipe_ready) begin
        counterValidAddrThreeStream_rValid <= 1'b0;
      end
      if(counterValidAddrThreeStream_s2mPipe_ready) begin
        counterValidAddrThreeStream_s2mPipe_rValid <= counterValidAddrThreeStream_s2mPipe_valid;
      end
      if(CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(counterValidAddrThreeStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_2 <= counterValidAddrThreeStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_12) begin
        CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_12) begin
        CICC1851_readStage_counterThreeValidStream_valid <= (CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready || CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_3);
      end
      if(controlStream_valid) begin
        controlStream_rValid <= 1'b1;
      end
      if(controlStream_s2mPipe_ready) begin
        controlStream_rValid <= 1'b0;
      end
      if(controlStream_s2mPipe_ready) begin
        controlStream_s2mPipe_rValid <= controlStream_s2mPipe_valid;
      end
      if(controlStream_s2mPipe_m2sPipe_ready) begin
        controlStream_s2mPipe_m2sPipe_rValid <= controlStream_s2mPipe_m2sPipe_valid;
      end
      if(controlStream_s2mPipe_m2sPipe_m2sPipe_valid) begin
        controlStream_s2mPipe_m2sPipe_m2sPipe_rValid <= 1'b1;
      end
      if(controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready) begin
        controlStream_s2mPipe_m2sPipe_m2sPipe_rValid <= 1'b0;
      end
      if(controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready) begin
        controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_valid;
      end
      if(readStage_mainOnePixelStream_valid) begin
        readStage_mainOnePixelStream_rValid <= 1'b1;
      end
      if(readStage_mainOnePixelStream_s2mPipe_ready) begin
        readStage_mainOnePixelStream_rValid <= 1'b0;
      end
      if(readStage_mainOnePixelStream_s2mPipe_ready) begin
        readStage_mainOnePixelStream_s2mPipe_rValid <= readStage_mainOnePixelStream_s2mPipe_valid;
      end
      if(readStage_counterOnePixelStream_valid) begin
        readStage_counterOnePixelStream_rValid <= 1'b1;
      end
      if(readStage_counterOnePixelStream_s2mPipe_ready) begin
        readStage_counterOnePixelStream_rValid <= 1'b0;
      end
      if(readStage_counterOnePixelStream_s2mPipe_ready) begin
        readStage_counterOnePixelStream_s2mPipe_rValid <= readStage_counterOnePixelStream_s2mPipe_valid;
      end
      if(readStage_mainTwoPixelStream_valid) begin
        readStage_mainTwoPixelStream_rValid <= 1'b1;
      end
      if(readStage_mainTwoPixelStream_s2mPipe_ready) begin
        readStage_mainTwoPixelStream_rValid <= 1'b0;
      end
      if(readStage_mainTwoPixelStream_s2mPipe_ready) begin
        readStage_mainTwoPixelStream_s2mPipe_rValid <= readStage_mainTwoPixelStream_s2mPipe_valid;
      end
      if(readStage_counterTwoPixelStream_valid) begin
        readStage_counterTwoPixelStream_rValid <= 1'b1;
      end
      if(readStage_counterTwoPixelStream_s2mPipe_ready) begin
        readStage_counterTwoPixelStream_rValid <= 1'b0;
      end
      if(readStage_counterTwoPixelStream_s2mPipe_ready) begin
        readStage_counterTwoPixelStream_s2mPipe_rValid <= readStage_counterTwoPixelStream_s2mPipe_valid;
      end
      if(readStage_mainThreePixelStream_valid) begin
        readStage_mainThreePixelStream_rValid <= 1'b1;
      end
      if(readStage_mainThreePixelStream_s2mPipe_ready) begin
        readStage_mainThreePixelStream_rValid <= 1'b0;
      end
      if(readStage_mainThreePixelStream_s2mPipe_ready) begin
        readStage_mainThreePixelStream_s2mPipe_rValid <= readStage_mainThreePixelStream_s2mPipe_valid;
      end
      if(readStage_counterThreePixelStream_valid) begin
        readStage_counterThreePixelStream_rValid <= 1'b1;
      end
      if(readStage_counterThreePixelStream_s2mPipe_ready) begin
        readStage_counterThreePixelStream_rValid <= 1'b0;
      end
      if(readStage_counterThreePixelStream_s2mPipe_ready) begin
        readStage_counterThreePixelStream_s2mPipe_rValid <= readStage_counterThreePixelStream_s2mPipe_valid;
      end
      if(readStage_mainOneValidStream_valid) begin
        readStage_mainOneValidStream_rValid <= 1'b1;
      end
      if(readStage_mainOneValidStream_s2mPipe_ready) begin
        readStage_mainOneValidStream_rValid <= 1'b0;
      end
      if(readStage_mainOneValidStream_s2mPipe_ready) begin
        readStage_mainOneValidStream_s2mPipe_rValid <= readStage_mainOneValidStream_s2mPipe_valid;
      end
      if(readStage_counterOneValidStream_valid) begin
        readStage_counterOneValidStream_rValid <= 1'b1;
      end
      if(readStage_counterOneValidStream_s2mPipe_ready) begin
        readStage_counterOneValidStream_rValid <= 1'b0;
      end
      if(readStage_counterOneValidStream_s2mPipe_ready) begin
        readStage_counterOneValidStream_s2mPipe_rValid <= readStage_counterOneValidStream_s2mPipe_valid;
      end
      if(readStage_mainTwoValidStream_valid) begin
        readStage_mainTwoValidStream_rValid <= 1'b1;
      end
      if(readStage_mainTwoValidStream_s2mPipe_ready) begin
        readStage_mainTwoValidStream_rValid <= 1'b0;
      end
      if(readStage_mainTwoValidStream_s2mPipe_ready) begin
        readStage_mainTwoValidStream_s2mPipe_rValid <= readStage_mainTwoValidStream_s2mPipe_valid;
      end
      if(readStage_counterTwoValidStream_valid) begin
        readStage_counterTwoValidStream_rValid <= 1'b1;
      end
      if(readStage_counterTwoValidStream_s2mPipe_ready) begin
        readStage_counterTwoValidStream_rValid <= 1'b0;
      end
      if(readStage_counterTwoValidStream_s2mPipe_ready) begin
        readStage_counterTwoValidStream_s2mPipe_rValid <= readStage_counterTwoValidStream_s2mPipe_valid;
      end
      if(readStage_mainThreeValidStream_valid) begin
        readStage_mainThreeValidStream_rValid <= 1'b1;
      end
      if(readStage_mainThreeValidStream_s2mPipe_ready) begin
        readStage_mainThreeValidStream_rValid <= 1'b0;
      end
      if(readStage_mainThreeValidStream_s2mPipe_ready) begin
        readStage_mainThreeValidStream_s2mPipe_rValid <= readStage_mainThreeValidStream_s2mPipe_valid;
      end
      if(readStage_counterThreeValidStream_valid) begin
        readStage_counterThreeValidStream_rValid <= 1'b1;
      end
      if(readStage_counterThreeValidStream_s2mPipe_ready) begin
        readStage_counterThreeValidStream_rValid <= 1'b0;
      end
      if(readStage_counterThreeValidStream_s2mPipe_ready) begin
        readStage_counterThreeValidStream_s2mPipe_rValid <= readStage_counterThreeValidStream_s2mPipe_valid;
      end
      if(readStage_controlPipe_translated_valid) begin
        readStage_controlPipe_translated_rValid <= 1'b1;
      end
      if(readStage_controlPipe_translated_s2mPipe_ready) begin
        readStage_controlPipe_translated_rValid <= 1'b0;
      end
      if(readStage_controlPipe_translated_s2mPipe_ready) begin
        readStage_controlPipe_translated_s2mPipe_rValid <= readStage_controlPipe_translated_s2mPipe_valid;
      end
      if(compareStage_mainOnePixelStream_valid) begin
        compareStage_mainOnePixelStream_rValid <= 1'b1;
      end
      if(compareStage_mainOnePixelStream_s2mPipe_ready) begin
        compareStage_mainOnePixelStream_rValid <= 1'b0;
      end
      if(compareStage_mainOnePixelStream_s2mPipe_ready) begin
        compareStage_mainOnePixelStream_s2mPipe_rValid <= compareStage_mainOnePixelStream_s2mPipe_valid;
      end
      if(compareStage_counterOnePixelStream_valid) begin
        compareStage_counterOnePixelStream_rValid <= 1'b1;
      end
      if(compareStage_counterOnePixelStream_s2mPipe_ready) begin
        compareStage_counterOnePixelStream_rValid <= 1'b0;
      end
      if(compareStage_counterOnePixelStream_s2mPipe_ready) begin
        compareStage_counterOnePixelStream_s2mPipe_rValid <= compareStage_counterOnePixelStream_s2mPipe_valid;
      end
      if(compareStage_mainTwoPixelStream_valid) begin
        compareStage_mainTwoPixelStream_rValid <= 1'b1;
      end
      if(compareStage_mainTwoPixelStream_s2mPipe_ready) begin
        compareStage_mainTwoPixelStream_rValid <= 1'b0;
      end
      if(compareStage_mainTwoPixelStream_s2mPipe_ready) begin
        compareStage_mainTwoPixelStream_s2mPipe_rValid <= compareStage_mainTwoPixelStream_s2mPipe_valid;
      end
      if(compareStage_counterTwoPixelStream_valid) begin
        compareStage_counterTwoPixelStream_rValid <= 1'b1;
      end
      if(compareStage_counterTwoPixelStream_s2mPipe_ready) begin
        compareStage_counterTwoPixelStream_rValid <= 1'b0;
      end
      if(compareStage_counterTwoPixelStream_s2mPipe_ready) begin
        compareStage_counterTwoPixelStream_s2mPipe_rValid <= compareStage_counterTwoPixelStream_s2mPipe_valid;
      end
      if(compareStage_mainThreePixelStream_valid) begin
        compareStage_mainThreePixelStream_rValid <= 1'b1;
      end
      if(compareStage_mainThreePixelStream_s2mPipe_ready) begin
        compareStage_mainThreePixelStream_rValid <= 1'b0;
      end
      if(compareStage_mainThreePixelStream_s2mPipe_ready) begin
        compareStage_mainThreePixelStream_s2mPipe_rValid <= compareStage_mainThreePixelStream_s2mPipe_valid;
      end
      if(compareStage_counterThreePixelStream_valid) begin
        compareStage_counterThreePixelStream_rValid <= 1'b1;
      end
      if(compareStage_counterThreePixelStream_s2mPipe_ready) begin
        compareStage_counterThreePixelStream_rValid <= 1'b0;
      end
      if(compareStage_counterThreePixelStream_s2mPipe_ready) begin
        compareStage_counterThreePixelStream_s2mPipe_rValid <= compareStage_counterThreePixelStream_s2mPipe_valid;
      end
      if(compareStage_mainOneValidStream_valid) begin
        compareStage_mainOneValidStream_rValid <= 1'b1;
      end
      if(compareStage_mainOneValidStream_s2mPipe_ready) begin
        compareStage_mainOneValidStream_rValid <= 1'b0;
      end
      if(compareStage_mainOneValidStream_s2mPipe_ready) begin
        compareStage_mainOneValidStream_s2mPipe_rValid <= compareStage_mainOneValidStream_s2mPipe_valid;
      end
      if(compareStage_counterOneValidStream_valid) begin
        compareStage_counterOneValidStream_rValid <= 1'b1;
      end
      if(compareStage_counterOneValidStream_s2mPipe_ready) begin
        compareStage_counterOneValidStream_rValid <= 1'b0;
      end
      if(compareStage_counterOneValidStream_s2mPipe_ready) begin
        compareStage_counterOneValidStream_s2mPipe_rValid <= compareStage_counterOneValidStream_s2mPipe_valid;
      end
      if(compareStage_mainTwoValidStream_valid) begin
        compareStage_mainTwoValidStream_rValid <= 1'b1;
      end
      if(compareStage_mainTwoValidStream_s2mPipe_ready) begin
        compareStage_mainTwoValidStream_rValid <= 1'b0;
      end
      if(compareStage_mainTwoValidStream_s2mPipe_ready) begin
        compareStage_mainTwoValidStream_s2mPipe_rValid <= compareStage_mainTwoValidStream_s2mPipe_valid;
      end
      if(compareStage_counterTwoValidStream_valid) begin
        compareStage_counterTwoValidStream_rValid <= 1'b1;
      end
      if(compareStage_counterTwoValidStream_s2mPipe_ready) begin
        compareStage_counterTwoValidStream_rValid <= 1'b0;
      end
      if(compareStage_counterTwoValidStream_s2mPipe_ready) begin
        compareStage_counterTwoValidStream_s2mPipe_rValid <= compareStage_counterTwoValidStream_s2mPipe_valid;
      end
      if(compareStage_mainThreeValidStream_valid) begin
        compareStage_mainThreeValidStream_rValid <= 1'b1;
      end
      if(compareStage_mainThreeValidStream_s2mPipe_ready) begin
        compareStage_mainThreeValidStream_rValid <= 1'b0;
      end
      if(compareStage_mainThreeValidStream_s2mPipe_ready) begin
        compareStage_mainThreeValidStream_s2mPipe_rValid <= compareStage_mainThreeValidStream_s2mPipe_valid;
      end
      if(compareStage_counterThreeValidStream_valid) begin
        compareStage_counterThreeValidStream_rValid <= 1'b1;
      end
      if(compareStage_counterThreeValidStream_s2mPipe_ready) begin
        compareStage_counterThreeValidStream_rValid <= 1'b0;
      end
      if(compareStage_counterThreeValidStream_s2mPipe_ready) begin
        compareStage_counterThreeValidStream_s2mPipe_rValid <= compareStage_counterThreeValidStream_s2mPipe_valid;
      end
      if(compareStage_controlPipe_translated_valid) begin
        compareStage_controlPipe_translated_rValid <= 1'b1;
      end
      if(compareStage_controlPipe_translated_s2mPipe_ready) begin
        compareStage_controlPipe_translated_rValid <= 1'b0;
      end
      if(compareStage_controlPipe_translated_s2mPipe_ready) begin
        compareStage_controlPipe_translated_s2mPipe_rValid <= compareStage_controlPipe_translated_s2mPipe_valid;
      end
      if(diffStage_mainOnePixelStream_valid) begin
        diffStage_mainOnePixelStream_rValid <= 1'b1;
      end
      if(diffStage_mainOnePixelStream_s2mPipe_ready) begin
        diffStage_mainOnePixelStream_rValid <= 1'b0;
      end
      if(diffStage_mainOnePixelStream_s2mPipe_ready) begin
        diffStage_mainOnePixelStream_s2mPipe_rValid <= diffStage_mainOnePixelStream_s2mPipe_valid;
      end
      if(diffStage_counterOnePixelStream_valid) begin
        diffStage_counterOnePixelStream_rValid <= 1'b1;
      end
      if(diffStage_counterOnePixelStream_s2mPipe_ready) begin
        diffStage_counterOnePixelStream_rValid <= 1'b0;
      end
      if(diffStage_counterOnePixelStream_s2mPipe_ready) begin
        diffStage_counterOnePixelStream_s2mPipe_rValid <= diffStage_counterOnePixelStream_s2mPipe_valid;
      end
      if(diffStage_mainTwoPixelStream_valid) begin
        diffStage_mainTwoPixelStream_rValid <= 1'b1;
      end
      if(diffStage_mainTwoPixelStream_s2mPipe_ready) begin
        diffStage_mainTwoPixelStream_rValid <= 1'b0;
      end
      if(diffStage_mainTwoPixelStream_s2mPipe_ready) begin
        diffStage_mainTwoPixelStream_s2mPipe_rValid <= diffStage_mainTwoPixelStream_s2mPipe_valid;
      end
      if(diffStage_counterTwoPixelStream_valid) begin
        diffStage_counterTwoPixelStream_rValid <= 1'b1;
      end
      if(diffStage_counterTwoPixelStream_s2mPipe_ready) begin
        diffStage_counterTwoPixelStream_rValid <= 1'b0;
      end
      if(diffStage_counterTwoPixelStream_s2mPipe_ready) begin
        diffStage_counterTwoPixelStream_s2mPipe_rValid <= diffStage_counterTwoPixelStream_s2mPipe_valid;
      end
      if(diffStage_mainThreePixelStream_valid) begin
        diffStage_mainThreePixelStream_rValid <= 1'b1;
      end
      if(diffStage_mainThreePixelStream_s2mPipe_ready) begin
        diffStage_mainThreePixelStream_rValid <= 1'b0;
      end
      if(diffStage_mainThreePixelStream_s2mPipe_ready) begin
        diffStage_mainThreePixelStream_s2mPipe_rValid <= diffStage_mainThreePixelStream_s2mPipe_valid;
      end
      if(diffStage_counterThreePixelStream_valid) begin
        diffStage_counterThreePixelStream_rValid <= 1'b1;
      end
      if(diffStage_counterThreePixelStream_s2mPipe_ready) begin
        diffStage_counterThreePixelStream_rValid <= 1'b0;
      end
      if(diffStage_counterThreePixelStream_s2mPipe_ready) begin
        diffStage_counterThreePixelStream_s2mPipe_rValid <= diffStage_counterThreePixelStream_s2mPipe_valid;
      end
      if(diffStage_mainOneValidStream_valid) begin
        diffStage_mainOneValidStream_rValid <= 1'b1;
      end
      if(diffStage_mainOneValidStream_s2mPipe_ready) begin
        diffStage_mainOneValidStream_rValid <= 1'b0;
      end
      if(diffStage_mainOneValidStream_s2mPipe_ready) begin
        diffStage_mainOneValidStream_s2mPipe_rValid <= diffStage_mainOneValidStream_s2mPipe_valid;
      end
      if(diffStage_counterOneValidStream_valid) begin
        diffStage_counterOneValidStream_rValid <= 1'b1;
      end
      if(diffStage_counterOneValidStream_s2mPipe_ready) begin
        diffStage_counterOneValidStream_rValid <= 1'b0;
      end
      if(diffStage_counterOneValidStream_s2mPipe_ready) begin
        diffStage_counterOneValidStream_s2mPipe_rValid <= diffStage_counterOneValidStream_s2mPipe_valid;
      end
      if(diffStage_mainTwoValidStream_valid) begin
        diffStage_mainTwoValidStream_rValid <= 1'b1;
      end
      if(diffStage_mainTwoValidStream_s2mPipe_ready) begin
        diffStage_mainTwoValidStream_rValid <= 1'b0;
      end
      if(diffStage_mainTwoValidStream_s2mPipe_ready) begin
        diffStage_mainTwoValidStream_s2mPipe_rValid <= diffStage_mainTwoValidStream_s2mPipe_valid;
      end
      if(diffStage_counterTwoValidStream_valid) begin
        diffStage_counterTwoValidStream_rValid <= 1'b1;
      end
      if(diffStage_counterTwoValidStream_s2mPipe_ready) begin
        diffStage_counterTwoValidStream_rValid <= 1'b0;
      end
      if(diffStage_counterTwoValidStream_s2mPipe_ready) begin
        diffStage_counterTwoValidStream_s2mPipe_rValid <= diffStage_counterTwoValidStream_s2mPipe_valid;
      end
      if(diffStage_mainThreeValidStream_valid) begin
        diffStage_mainThreeValidStream_rValid <= 1'b1;
      end
      if(diffStage_mainThreeValidStream_s2mPipe_ready) begin
        diffStage_mainThreeValidStream_rValid <= 1'b0;
      end
      if(diffStage_mainThreeValidStream_s2mPipe_ready) begin
        diffStage_mainThreeValidStream_s2mPipe_rValid <= diffStage_mainThreeValidStream_s2mPipe_valid;
      end
      if(diffStage_counterThreeValidStream_valid) begin
        diffStage_counterThreeValidStream_rValid <= 1'b1;
      end
      if(diffStage_counterThreeValidStream_s2mPipe_ready) begin
        diffStage_counterThreeValidStream_rValid <= 1'b0;
      end
      if(diffStage_counterThreeValidStream_s2mPipe_ready) begin
        diffStage_counterThreeValidStream_s2mPipe_rValid <= diffStage_counterThreeValidStream_s2mPipe_valid;
      end
      if(resultStage_controlPipeBeforePipe_valid) begin
        resultStage_controlPipeBeforePipe_rValid <= 1'b1;
      end
      if(resultStage_controlPipeBeforePipe_s2mPipe_ready) begin
        resultStage_controlPipeBeforePipe_rValid <= 1'b0;
      end
      if(resultStage_controlPipeBeforePipe_s2mPipe_ready) begin
        resultStage_controlPipeBeforePipe_s2mPipe_rValid <= resultStage_controlPipeBeforePipe_s2mPipe_valid;
      end
      if(resultStage_pixelStream_valid) begin
        resultStage_pixelStream_rValid <= 1'b1;
      end
      if(resultStage_pixelStream_s2mPipe_ready) begin
        resultStage_pixelStream_rValid <= 1'b0;
      end
      if(resultStage_pixelStream_s2mPipe_ready) begin
        resultStage_pixelStream_s2mPipe_rValid <= resultStage_pixelStream_s2mPipe_valid;
      end
      if(when_SuperResolutionPart3_l1115) begin
        isHorizontalDirection <= resultStage_controlPipeBeforePipe_payload_isHorizontalMin;
        minDiff <= resultStage_controlPipeBeforePipe_payload_minDiff;
        candidatePixel <= resultStage_pixelStream_payload;
      end
      if(diffStage_controlPipe_fire) begin
        inValidMinDiff <= diffStage_controlPipe_payload_inValidMinDiff;
      end
      if(pixelsStream_valid) begin
        pixelsStream_rValid <= 1'b1;
      end
      if(pixelsStream_s2mPipe_ready) begin
        pixelsStream_rValid <= 1'b0;
      end
      if(pixelsStream_s2mPipe_ready) begin
        pixelsStream_s2mPipe_rValid <= pixelsStream_s2mPipe_valid;
      end
      controlStateMachine_stateReg <= controlStateMachine_stateNext;
      case(controlStateMachine_stateReg)
        controlStateMachine_enumDef_8_HOLD : begin
        end
        controlStateMachine_enumDef_8_PASS : begin
        end
        controlStateMachine_enumDef_8_EXTRA : begin
          if(when_SuperResolutionPart3_l1220) begin
            frameStart <= 1'b0;
          end
          if(when_SuperResolutionPart3_l1223) begin
            outReachRowEnd <= 1'b1;
          end
          if(when_SuperResolutionPart3_l1224) begin
            outReachFinalRow <= 1'b1;
          end
          if(when_SuperResolutionPart3_l1226) begin
            if(outReachFinalRow) begin
              startRead <= 1'b0;
              readDone <= 1'b1;
              outReachRowEnd <= 1'b0;
              outReachFinalRow <= 1'b0;
            end else begin
              outReachRowEnd <= 1'b0;
            end
          end
          if(controlStream_fire_6) begin
            if(outReachRowEnd) begin
              outReachRowEnd <= 1'b0;
            end
          end
          if(when_SuperResolutionPart3_l1247) begin
            if(when_SuperResolutionPart3_l1248) begin
              holdBuffer <= 1'b0;
            end
            if(when_SuperResolutionPart3_l1250) begin
              currentRowBuffer <= 2'b00;
            end else begin
              currentRowBuffer <= (currentRowBuffer + 2'b01);
            end
            if(when_SuperResolutionPart3_l1252) begin
              nextRowBuffer <= 2'b00;
            end else begin
              nextRowBuffer <= (nextRowBuffer + 2'b01);
            end
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(posedge clk) begin
    startIn_regNext <= startIn;
    startIn_regNext_1 <= startIn;
    if(pixelsIn_ready) begin
      pixelsIn_rData_pixel <= pixelsIn_payload_pixel;
      pixelsIn_rData_frameStart <= pixelsIn_payload_frameStart;
      pixelsIn_rData_rowEnd <= pixelsIn_payload_rowEnd;
      pixelsIn_rData_inpValid <= pixelsIn_payload_inpValid;
    end
    if(pixelsIn_s2mPipe_ready) begin
      pixelsIn_s2mPipe_rData_pixel <= pixelsIn_s2mPipe_payload_pixel;
      pixelsIn_s2mPipe_rData_frameStart <= pixelsIn_s2mPipe_payload_frameStart;
      pixelsIn_s2mPipe_rData_rowEnd <= pixelsIn_s2mPipe_payload_rowEnd;
      pixelsIn_s2mPipe_rData_inpValid <= pixelsIn_s2mPipe_payload_inpValid;
    end
    if(mainPixelAddrOneStream_ready) begin
      mainPixelAddrOneStream_rData <= mainPixelAddrOneStream_payload;
    end
    if(mainPixelAddrOneStream_s2mPipe_ready) begin
      mainPixelAddrOneStream_s2mPipe_rData <= mainPixelAddrOneStream_s2mPipe_payload;
    end
    if(CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_mainOnePixelStream_payload_1 <= CICC1851_readStage_mainOnePixelStream_payload;
    end
    if(CICC1851_1) begin
      CICC1851_readStage_mainOnePixelStream_payload_2 <= (CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_mainOnePixelStream_payload_1 : CICC1851_readStage_mainOnePixelStream_payload);
    end
    if(counterPixelAddrOneStream_ready) begin
      counterPixelAddrOneStream_rData <= counterPixelAddrOneStream_payload;
    end
    if(counterPixelAddrOneStream_s2mPipe_ready) begin
      counterPixelAddrOneStream_s2mPipe_rData <= counterPixelAddrOneStream_s2mPipe_payload;
    end
    if(CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_counterOnePixelStream_payload_1 <= CICC1851_readStage_counterOnePixelStream_payload;
    end
    if(CICC1851_2) begin
      CICC1851_readStage_counterOnePixelStream_payload_2 <= (CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_counterOnePixelStream_payload_1 : CICC1851_readStage_counterOnePixelStream_payload);
    end
    if(mainPixelAddrTwoStream_ready) begin
      mainPixelAddrTwoStream_rData <= mainPixelAddrTwoStream_payload;
    end
    if(mainPixelAddrTwoStream_s2mPipe_ready) begin
      mainPixelAddrTwoStream_s2mPipe_rData <= mainPixelAddrTwoStream_s2mPipe_payload;
    end
    if(CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_mainTwoPixelStream_payload_1 <= CICC1851_readStage_mainTwoPixelStream_payload;
    end
    if(CICC1851_3) begin
      CICC1851_readStage_mainTwoPixelStream_payload_2 <= (CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_mainTwoPixelStream_payload_1 : CICC1851_readStage_mainTwoPixelStream_payload);
    end
    if(counterPixelAddrTwoStream_ready) begin
      counterPixelAddrTwoStream_rData <= counterPixelAddrTwoStream_payload;
    end
    if(counterPixelAddrTwoStream_s2mPipe_ready) begin
      counterPixelAddrTwoStream_s2mPipe_rData <= counterPixelAddrTwoStream_s2mPipe_payload;
    end
    if(CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_counterTwoPixelStream_payload_1 <= CICC1851_readStage_counterTwoPixelStream_payload;
    end
    if(CICC1851_4) begin
      CICC1851_readStage_counterTwoPixelStream_payload_2 <= (CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_counterTwoPixelStream_payload_1 : CICC1851_readStage_counterTwoPixelStream_payload);
    end
    if(mainPixelAddrThreeStream_ready) begin
      mainPixelAddrThreeStream_rData <= mainPixelAddrThreeStream_payload;
    end
    if(mainPixelAddrThreeStream_s2mPipe_ready) begin
      mainPixelAddrThreeStream_s2mPipe_rData <= mainPixelAddrThreeStream_s2mPipe_payload;
    end
    if(CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_mainThreePixelStream_payload_1 <= CICC1851_readStage_mainThreePixelStream_payload;
    end
    if(CICC1851_5) begin
      CICC1851_readStage_mainThreePixelStream_payload_2 <= (CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_mainThreePixelStream_payload_1 : CICC1851_readStage_mainThreePixelStream_payload);
    end
    if(counterPixelAddrThreeStream_ready) begin
      counterPixelAddrThreeStream_rData <= counterPixelAddrThreeStream_payload;
    end
    if(counterPixelAddrThreeStream_s2mPipe_ready) begin
      counterPixelAddrThreeStream_s2mPipe_rData <= counterPixelAddrThreeStream_s2mPipe_payload;
    end
    if(CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_counterThreePixelStream_payload_1 <= CICC1851_readStage_counterThreePixelStream_payload;
    end
    if(CICC1851_6) begin
      CICC1851_readStage_counterThreePixelStream_payload_2 <= (CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_counterThreePixelStream_payload_1 : CICC1851_readStage_counterThreePixelStream_payload);
    end
    if(mainValidAddrOneStream_ready) begin
      mainValidAddrOneStream_rData <= mainValidAddrOneStream_payload;
    end
    if(mainValidAddrOneStream_s2mPipe_ready) begin
      mainValidAddrOneStream_s2mPipe_rData <= mainValidAddrOneStream_s2mPipe_payload;
    end
    if(CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_mainOneValidStream_payload_1 <= CICC1851_readStage_mainOneValidStream_payload;
    end
    if(CICC1851_7) begin
      CICC1851_readStage_mainOneValidStream_payload_2 <= (CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_mainOneValidStream_payload_1 : CICC1851_readStage_mainOneValidStream_payload);
    end
    if(counterValidAddrOneStream_ready) begin
      counterValidAddrOneStream_rData <= counterValidAddrOneStream_payload;
    end
    if(counterValidAddrOneStream_s2mPipe_ready) begin
      counterValidAddrOneStream_s2mPipe_rData <= counterValidAddrOneStream_s2mPipe_payload;
    end
    if(CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_counterOneValidStream_payload_1 <= CICC1851_readStage_counterOneValidStream_payload;
    end
    if(CICC1851_8) begin
      CICC1851_readStage_counterOneValidStream_payload_2 <= (CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_counterOneValidStream_payload_1 : CICC1851_readStage_counterOneValidStream_payload);
    end
    if(mainValidAddrTwoStream_ready) begin
      mainValidAddrTwoStream_rData <= mainValidAddrTwoStream_payload;
    end
    if(mainValidAddrTwoStream_s2mPipe_ready) begin
      mainValidAddrTwoStream_s2mPipe_rData <= mainValidAddrTwoStream_s2mPipe_payload;
    end
    if(CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_mainTwoValidStream_payload_1 <= CICC1851_readStage_mainTwoValidStream_payload;
    end
    if(CICC1851_9) begin
      CICC1851_readStage_mainTwoValidStream_payload_2 <= (CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_mainTwoValidStream_payload_1 : CICC1851_readStage_mainTwoValidStream_payload);
    end
    if(counterValidAddrTwoStream_ready) begin
      counterValidAddrTwoStream_rData <= counterValidAddrTwoStream_payload;
    end
    if(counterValidAddrTwoStream_s2mPipe_ready) begin
      counterValidAddrTwoStream_s2mPipe_rData <= counterValidAddrTwoStream_s2mPipe_payload;
    end
    if(CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_counterTwoValidStream_payload_1 <= CICC1851_readStage_counterTwoValidStream_payload;
    end
    if(CICC1851_10) begin
      CICC1851_readStage_counterTwoValidStream_payload_2 <= (CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_counterTwoValidStream_payload_1 : CICC1851_readStage_counterTwoValidStream_payload);
    end
    if(mainValidAddrThreeStream_ready) begin
      mainValidAddrThreeStream_rData <= mainValidAddrThreeStream_payload;
    end
    if(mainValidAddrThreeStream_s2mPipe_ready) begin
      mainValidAddrThreeStream_s2mPipe_rData <= mainValidAddrThreeStream_s2mPipe_payload;
    end
    if(CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_mainThreeValidStream_payload_1 <= CICC1851_readStage_mainThreeValidStream_payload;
    end
    if(CICC1851_11) begin
      CICC1851_readStage_mainThreeValidStream_payload_2 <= (CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_mainThreeValidStream_payload_1 : CICC1851_readStage_mainThreeValidStream_payload);
    end
    if(counterValidAddrThreeStream_ready) begin
      counterValidAddrThreeStream_rData <= counterValidAddrThreeStream_payload;
    end
    if(counterValidAddrThreeStream_s2mPipe_ready) begin
      counterValidAddrThreeStream_s2mPipe_rData <= counterValidAddrThreeStream_s2mPipe_payload;
    end
    if(CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_counterThreeValidStream_payload_1 <= CICC1851_readStage_counterThreeValidStream_payload;
    end
    if(CICC1851_12) begin
      CICC1851_readStage_counterThreeValidStream_payload_2 <= (CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_counterThreeValidStream_payload_1 : CICC1851_readStage_counterThreeValidStream_payload);
    end
    if(controlStream_ready) begin
      controlStream_rData_frameStart <= controlStream_payload_frameStart;
      controlStream_rData_rowEnd <= controlStream_payload_rowEnd;
      controlStream_rData_pipeValid <= controlStream_payload_pipeValid;
      controlStream_rData_firstRow <= controlStream_payload_firstRow;
      controlStream_rData_lastRow <= controlStream_payload_lastRow;
      controlStream_rData_finalResult <= controlStream_payload_finalResult;
      controlStream_rData_mainCompare <= controlStream_payload_mainCompare;
      controlStream_rData_counterCompare <= controlStream_payload_counterCompare;
      controlStream_rData_horizontalCompare <= controlStream_payload_horizontalCompare;
      controlStream_rData_verticalCompare <= controlStream_payload_verticalCompare;
      controlStream_rData_mainDiff <= controlStream_payload_mainDiff;
      controlStream_rData_counterDiff <= controlStream_payload_counterDiff;
      controlStream_rData_horizontalDiff <= controlStream_payload_horizontalDiff;
      controlStream_rData_verticalDiff <= controlStream_payload_verticalDiff;
      controlStream_rData_isHorizontalMin <= controlStream_payload_isHorizontalMin;
      controlStream_rData_minDiff <= controlStream_payload_minDiff;
      controlStream_rData_currentPosition <= controlStream_payload_currentPosition;
      controlStream_rData_nextPosition <= controlStream_payload_nextPosition;
      controlStream_rData_horizontalDirectionValid <= controlStream_payload_horizontalDirectionValid;
      controlStream_rData_verticalDirectionValid <= controlStream_payload_verticalDirectionValid;
      controlStream_rData_mainDirectionValid <= controlStream_payload_mainDirectionValid;
      controlStream_rData_counterDirectionValid <= controlStream_payload_counterDirectionValid;
      controlStream_rData_inValidMinDiff <= controlStream_payload_inValidMinDiff;
    end
    if(controlStream_s2mPipe_ready) begin
      controlStream_s2mPipe_rData_frameStart <= controlStream_s2mPipe_payload_frameStart;
      controlStream_s2mPipe_rData_rowEnd <= controlStream_s2mPipe_payload_rowEnd;
      controlStream_s2mPipe_rData_pipeValid <= controlStream_s2mPipe_payload_pipeValid;
      controlStream_s2mPipe_rData_firstRow <= controlStream_s2mPipe_payload_firstRow;
      controlStream_s2mPipe_rData_lastRow <= controlStream_s2mPipe_payload_lastRow;
      controlStream_s2mPipe_rData_finalResult <= controlStream_s2mPipe_payload_finalResult;
      controlStream_s2mPipe_rData_mainCompare <= controlStream_s2mPipe_payload_mainCompare;
      controlStream_s2mPipe_rData_counterCompare <= controlStream_s2mPipe_payload_counterCompare;
      controlStream_s2mPipe_rData_horizontalCompare <= controlStream_s2mPipe_payload_horizontalCompare;
      controlStream_s2mPipe_rData_verticalCompare <= controlStream_s2mPipe_payload_verticalCompare;
      controlStream_s2mPipe_rData_mainDiff <= controlStream_s2mPipe_payload_mainDiff;
      controlStream_s2mPipe_rData_counterDiff <= controlStream_s2mPipe_payload_counterDiff;
      controlStream_s2mPipe_rData_horizontalDiff <= controlStream_s2mPipe_payload_horizontalDiff;
      controlStream_s2mPipe_rData_verticalDiff <= controlStream_s2mPipe_payload_verticalDiff;
      controlStream_s2mPipe_rData_isHorizontalMin <= controlStream_s2mPipe_payload_isHorizontalMin;
      controlStream_s2mPipe_rData_minDiff <= controlStream_s2mPipe_payload_minDiff;
      controlStream_s2mPipe_rData_currentPosition <= controlStream_s2mPipe_payload_currentPosition;
      controlStream_s2mPipe_rData_nextPosition <= controlStream_s2mPipe_payload_nextPosition;
      controlStream_s2mPipe_rData_horizontalDirectionValid <= controlStream_s2mPipe_payload_horizontalDirectionValid;
      controlStream_s2mPipe_rData_verticalDirectionValid <= controlStream_s2mPipe_payload_verticalDirectionValid;
      controlStream_s2mPipe_rData_mainDirectionValid <= controlStream_s2mPipe_payload_mainDirectionValid;
      controlStream_s2mPipe_rData_counterDirectionValid <= controlStream_s2mPipe_payload_counterDirectionValid;
      controlStream_s2mPipe_rData_inValidMinDiff <= controlStream_s2mPipe_payload_inValidMinDiff;
    end
    if(controlStream_s2mPipe_m2sPipe_ready) begin
      controlStream_s2mPipe_m2sPipe_rData_frameStart <= controlStream_s2mPipe_m2sPipe_payload_frameStart;
      controlStream_s2mPipe_m2sPipe_rData_rowEnd <= controlStream_s2mPipe_m2sPipe_payload_rowEnd;
      controlStream_s2mPipe_m2sPipe_rData_pipeValid <= controlStream_s2mPipe_m2sPipe_payload_pipeValid;
      controlStream_s2mPipe_m2sPipe_rData_firstRow <= controlStream_s2mPipe_m2sPipe_payload_firstRow;
      controlStream_s2mPipe_m2sPipe_rData_lastRow <= controlStream_s2mPipe_m2sPipe_payload_lastRow;
      controlStream_s2mPipe_m2sPipe_rData_finalResult <= controlStream_s2mPipe_m2sPipe_payload_finalResult;
      controlStream_s2mPipe_m2sPipe_rData_mainCompare <= controlStream_s2mPipe_m2sPipe_payload_mainCompare;
      controlStream_s2mPipe_m2sPipe_rData_counterCompare <= controlStream_s2mPipe_m2sPipe_payload_counterCompare;
      controlStream_s2mPipe_m2sPipe_rData_horizontalCompare <= controlStream_s2mPipe_m2sPipe_payload_horizontalCompare;
      controlStream_s2mPipe_m2sPipe_rData_verticalCompare <= controlStream_s2mPipe_m2sPipe_payload_verticalCompare;
      controlStream_s2mPipe_m2sPipe_rData_mainDiff <= controlStream_s2mPipe_m2sPipe_payload_mainDiff;
      controlStream_s2mPipe_m2sPipe_rData_counterDiff <= controlStream_s2mPipe_m2sPipe_payload_counterDiff;
      controlStream_s2mPipe_m2sPipe_rData_horizontalDiff <= controlStream_s2mPipe_m2sPipe_payload_horizontalDiff;
      controlStream_s2mPipe_m2sPipe_rData_verticalDiff <= controlStream_s2mPipe_m2sPipe_payload_verticalDiff;
      controlStream_s2mPipe_m2sPipe_rData_isHorizontalMin <= controlStream_s2mPipe_m2sPipe_payload_isHorizontalMin;
      controlStream_s2mPipe_m2sPipe_rData_minDiff <= controlStream_s2mPipe_m2sPipe_payload_minDiff;
      controlStream_s2mPipe_m2sPipe_rData_currentPosition <= controlStream_s2mPipe_m2sPipe_payload_currentPosition;
      controlStream_s2mPipe_m2sPipe_rData_nextPosition <= controlStream_s2mPipe_m2sPipe_payload_nextPosition;
      controlStream_s2mPipe_m2sPipe_rData_horizontalDirectionValid <= controlStream_s2mPipe_m2sPipe_payload_horizontalDirectionValid;
      controlStream_s2mPipe_m2sPipe_rData_verticalDirectionValid <= controlStream_s2mPipe_m2sPipe_payload_verticalDirectionValid;
      controlStream_s2mPipe_m2sPipe_rData_mainDirectionValid <= controlStream_s2mPipe_m2sPipe_payload_mainDirectionValid;
      controlStream_s2mPipe_m2sPipe_rData_counterDirectionValid <= controlStream_s2mPipe_m2sPipe_payload_counterDirectionValid;
      controlStream_s2mPipe_m2sPipe_rData_inValidMinDiff <= controlStream_s2mPipe_m2sPipe_payload_inValidMinDiff;
    end
    if(controlStream_s2mPipe_m2sPipe_m2sPipe_ready) begin
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_frameStart <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_frameStart;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_rowEnd <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_rowEnd;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_pipeValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_pipeValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_firstRow <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_firstRow;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_lastRow <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_lastRow;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_finalResult <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_finalResult;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_horizontalCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_horizontalCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_verticalCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_verticalCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_horizontalDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_horizontalDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_verticalDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_verticalDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_isHorizontalMin <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_isHorizontalMin;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_minDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_minDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_currentPosition <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_currentPosition;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_nextPosition <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_nextPosition;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_horizontalDirectionValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_horizontalDirectionValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_verticalDirectionValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_verticalDirectionValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainDirectionValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDirectionValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterDirectionValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDirectionValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_inValidMinDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_inValidMinDiff;
    end
    if(controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready) begin
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_frameStart <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_frameStart;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_rowEnd <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_rowEnd;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_pipeValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_pipeValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_firstRow <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_firstRow;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_lastRow <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_lastRow;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_finalResult <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_finalResult;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_horizontalCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_horizontalCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_verticalCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_verticalCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_horizontalDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_horizontalDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_verticalDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_verticalDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_isHorizontalMin <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_isHorizontalMin;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_minDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_minDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_currentPosition <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_currentPosition;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_nextPosition <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_nextPosition;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_horizontalDirectionValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_horizontalDirectionValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_verticalDirectionValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_verticalDirectionValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainDirectionValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainDirectionValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterDirectionValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterDirectionValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_inValidMinDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_inValidMinDiff;
    end
    if(readStage_mainOnePixelStream_ready) begin
      readStage_mainOnePixelStream_rData <= readStage_mainOnePixelStream_payload;
    end
    if(readStage_mainOnePixelStream_s2mPipe_ready) begin
      readStage_mainOnePixelStream_s2mPipe_rData <= readStage_mainOnePixelStream_s2mPipe_payload;
    end
    if(readStage_counterOnePixelStream_ready) begin
      readStage_counterOnePixelStream_rData <= readStage_counterOnePixelStream_payload;
    end
    if(readStage_counterOnePixelStream_s2mPipe_ready) begin
      readStage_counterOnePixelStream_s2mPipe_rData <= readStage_counterOnePixelStream_s2mPipe_payload;
    end
    if(readStage_mainTwoPixelStream_ready) begin
      readStage_mainTwoPixelStream_rData <= readStage_mainTwoPixelStream_payload;
    end
    if(readStage_mainTwoPixelStream_s2mPipe_ready) begin
      readStage_mainTwoPixelStream_s2mPipe_rData <= readStage_mainTwoPixelStream_s2mPipe_payload;
    end
    if(readStage_counterTwoPixelStream_ready) begin
      readStage_counterTwoPixelStream_rData <= readStage_counterTwoPixelStream_payload;
    end
    if(readStage_counterTwoPixelStream_s2mPipe_ready) begin
      readStage_counterTwoPixelStream_s2mPipe_rData <= readStage_counterTwoPixelStream_s2mPipe_payload;
    end
    if(readStage_mainThreePixelStream_ready) begin
      readStage_mainThreePixelStream_rData <= readStage_mainThreePixelStream_payload;
    end
    if(readStage_mainThreePixelStream_s2mPipe_ready) begin
      readStage_mainThreePixelStream_s2mPipe_rData <= readStage_mainThreePixelStream_s2mPipe_payload;
    end
    if(readStage_counterThreePixelStream_ready) begin
      readStage_counterThreePixelStream_rData <= readStage_counterThreePixelStream_payload;
    end
    if(readStage_counterThreePixelStream_s2mPipe_ready) begin
      readStage_counterThreePixelStream_s2mPipe_rData <= readStage_counterThreePixelStream_s2mPipe_payload;
    end
    if(readStage_mainOneValidStream_ready) begin
      readStage_mainOneValidStream_rData <= readStage_mainOneValidStream_payload;
    end
    if(readStage_mainOneValidStream_s2mPipe_ready) begin
      readStage_mainOneValidStream_s2mPipe_rData <= readStage_mainOneValidStream_s2mPipe_payload;
    end
    if(readStage_counterOneValidStream_ready) begin
      readStage_counterOneValidStream_rData <= readStage_counterOneValidStream_payload;
    end
    if(readStage_counterOneValidStream_s2mPipe_ready) begin
      readStage_counterOneValidStream_s2mPipe_rData <= readStage_counterOneValidStream_s2mPipe_payload;
    end
    if(readStage_mainTwoValidStream_ready) begin
      readStage_mainTwoValidStream_rData <= readStage_mainTwoValidStream_payload;
    end
    if(readStage_mainTwoValidStream_s2mPipe_ready) begin
      readStage_mainTwoValidStream_s2mPipe_rData <= readStage_mainTwoValidStream_s2mPipe_payload;
    end
    if(readStage_counterTwoValidStream_ready) begin
      readStage_counterTwoValidStream_rData <= readStage_counterTwoValidStream_payload;
    end
    if(readStage_counterTwoValidStream_s2mPipe_ready) begin
      readStage_counterTwoValidStream_s2mPipe_rData <= readStage_counterTwoValidStream_s2mPipe_payload;
    end
    if(readStage_mainThreeValidStream_ready) begin
      readStage_mainThreeValidStream_rData <= readStage_mainThreeValidStream_payload;
    end
    if(readStage_mainThreeValidStream_s2mPipe_ready) begin
      readStage_mainThreeValidStream_s2mPipe_rData <= readStage_mainThreeValidStream_s2mPipe_payload;
    end
    if(readStage_counterThreeValidStream_ready) begin
      readStage_counterThreeValidStream_rData <= readStage_counterThreeValidStream_payload;
    end
    if(readStage_counterThreeValidStream_s2mPipe_ready) begin
      readStage_counterThreeValidStream_s2mPipe_rData <= readStage_counterThreeValidStream_s2mPipe_payload;
    end
    if(readStage_controlPipe_translated_ready) begin
      readStage_controlPipe_translated_rData_frameStart <= readStage_controlPipe_translated_payload_frameStart;
      readStage_controlPipe_translated_rData_rowEnd <= readStage_controlPipe_translated_payload_rowEnd;
      readStage_controlPipe_translated_rData_pipeValid <= readStage_controlPipe_translated_payload_pipeValid;
      readStage_controlPipe_translated_rData_firstRow <= readStage_controlPipe_translated_payload_firstRow;
      readStage_controlPipe_translated_rData_lastRow <= readStage_controlPipe_translated_payload_lastRow;
      readStage_controlPipe_translated_rData_finalResult <= readStage_controlPipe_translated_payload_finalResult;
      readStage_controlPipe_translated_rData_mainCompare <= readStage_controlPipe_translated_payload_mainCompare;
      readStage_controlPipe_translated_rData_counterCompare <= readStage_controlPipe_translated_payload_counterCompare;
      readStage_controlPipe_translated_rData_horizontalCompare <= readStage_controlPipe_translated_payload_horizontalCompare;
      readStage_controlPipe_translated_rData_verticalCompare <= readStage_controlPipe_translated_payload_verticalCompare;
      readStage_controlPipe_translated_rData_mainDiff <= readStage_controlPipe_translated_payload_mainDiff;
      readStage_controlPipe_translated_rData_counterDiff <= readStage_controlPipe_translated_payload_counterDiff;
      readStage_controlPipe_translated_rData_horizontalDiff <= readStage_controlPipe_translated_payload_horizontalDiff;
      readStage_controlPipe_translated_rData_verticalDiff <= readStage_controlPipe_translated_payload_verticalDiff;
      readStage_controlPipe_translated_rData_isHorizontalMin <= readStage_controlPipe_translated_payload_isHorizontalMin;
      readStage_controlPipe_translated_rData_minDiff <= readStage_controlPipe_translated_payload_minDiff;
      readStage_controlPipe_translated_rData_currentPosition <= readStage_controlPipe_translated_payload_currentPosition;
      readStage_controlPipe_translated_rData_nextPosition <= readStage_controlPipe_translated_payload_nextPosition;
      readStage_controlPipe_translated_rData_horizontalDirectionValid <= readStage_controlPipe_translated_payload_horizontalDirectionValid;
      readStage_controlPipe_translated_rData_verticalDirectionValid <= readStage_controlPipe_translated_payload_verticalDirectionValid;
      readStage_controlPipe_translated_rData_mainDirectionValid <= readStage_controlPipe_translated_payload_mainDirectionValid;
      readStage_controlPipe_translated_rData_counterDirectionValid <= readStage_controlPipe_translated_payload_counterDirectionValid;
      readStage_controlPipe_translated_rData_inValidMinDiff <= readStage_controlPipe_translated_payload_inValidMinDiff;
    end
    if(readStage_controlPipe_translated_s2mPipe_ready) begin
      readStage_controlPipe_translated_s2mPipe_rData_frameStart <= readStage_controlPipe_translated_s2mPipe_payload_frameStart;
      readStage_controlPipe_translated_s2mPipe_rData_rowEnd <= readStage_controlPipe_translated_s2mPipe_payload_rowEnd;
      readStage_controlPipe_translated_s2mPipe_rData_pipeValid <= readStage_controlPipe_translated_s2mPipe_payload_pipeValid;
      readStage_controlPipe_translated_s2mPipe_rData_firstRow <= readStage_controlPipe_translated_s2mPipe_payload_firstRow;
      readStage_controlPipe_translated_s2mPipe_rData_lastRow <= readStage_controlPipe_translated_s2mPipe_payload_lastRow;
      readStage_controlPipe_translated_s2mPipe_rData_finalResult <= readStage_controlPipe_translated_s2mPipe_payload_finalResult;
      readStage_controlPipe_translated_s2mPipe_rData_mainCompare <= readStage_controlPipe_translated_s2mPipe_payload_mainCompare;
      readStage_controlPipe_translated_s2mPipe_rData_counterCompare <= readStage_controlPipe_translated_s2mPipe_payload_counterCompare;
      readStage_controlPipe_translated_s2mPipe_rData_horizontalCompare <= readStage_controlPipe_translated_s2mPipe_payload_horizontalCompare;
      readStage_controlPipe_translated_s2mPipe_rData_verticalCompare <= readStage_controlPipe_translated_s2mPipe_payload_verticalCompare;
      readStage_controlPipe_translated_s2mPipe_rData_mainDiff <= readStage_controlPipe_translated_s2mPipe_payload_mainDiff;
      readStage_controlPipe_translated_s2mPipe_rData_counterDiff <= readStage_controlPipe_translated_s2mPipe_payload_counterDiff;
      readStage_controlPipe_translated_s2mPipe_rData_horizontalDiff <= readStage_controlPipe_translated_s2mPipe_payload_horizontalDiff;
      readStage_controlPipe_translated_s2mPipe_rData_verticalDiff <= readStage_controlPipe_translated_s2mPipe_payload_verticalDiff;
      readStage_controlPipe_translated_s2mPipe_rData_isHorizontalMin <= readStage_controlPipe_translated_s2mPipe_payload_isHorizontalMin;
      readStage_controlPipe_translated_s2mPipe_rData_minDiff <= readStage_controlPipe_translated_s2mPipe_payload_minDiff;
      readStage_controlPipe_translated_s2mPipe_rData_currentPosition <= readStage_controlPipe_translated_s2mPipe_payload_currentPosition;
      readStage_controlPipe_translated_s2mPipe_rData_nextPosition <= readStage_controlPipe_translated_s2mPipe_payload_nextPosition;
      readStage_controlPipe_translated_s2mPipe_rData_horizontalDirectionValid <= readStage_controlPipe_translated_s2mPipe_payload_horizontalDirectionValid;
      readStage_controlPipe_translated_s2mPipe_rData_verticalDirectionValid <= readStage_controlPipe_translated_s2mPipe_payload_verticalDirectionValid;
      readStage_controlPipe_translated_s2mPipe_rData_mainDirectionValid <= readStage_controlPipe_translated_s2mPipe_payload_mainDirectionValid;
      readStage_controlPipe_translated_s2mPipe_rData_counterDirectionValid <= readStage_controlPipe_translated_s2mPipe_payload_counterDirectionValid;
      readStage_controlPipe_translated_s2mPipe_rData_inValidMinDiff <= readStage_controlPipe_translated_s2mPipe_payload_inValidMinDiff;
    end
    if(compareStage_mainOnePixelStream_ready) begin
      compareStage_mainOnePixelStream_rData <= compareStage_mainOnePixelStream_payload;
    end
    if(compareStage_mainOnePixelStream_s2mPipe_ready) begin
      compareStage_mainOnePixelStream_s2mPipe_rData <= compareStage_mainOnePixelStream_s2mPipe_payload;
    end
    if(compareStage_counterOnePixelStream_ready) begin
      compareStage_counterOnePixelStream_rData <= compareStage_counterOnePixelStream_payload;
    end
    if(compareStage_counterOnePixelStream_s2mPipe_ready) begin
      compareStage_counterOnePixelStream_s2mPipe_rData <= compareStage_counterOnePixelStream_s2mPipe_payload;
    end
    if(compareStage_mainTwoPixelStream_ready) begin
      compareStage_mainTwoPixelStream_rData <= compareStage_mainTwoPixelStream_payload;
    end
    if(compareStage_mainTwoPixelStream_s2mPipe_ready) begin
      compareStage_mainTwoPixelStream_s2mPipe_rData <= compareStage_mainTwoPixelStream_s2mPipe_payload;
    end
    if(compareStage_counterTwoPixelStream_ready) begin
      compareStage_counterTwoPixelStream_rData <= compareStage_counterTwoPixelStream_payload;
    end
    if(compareStage_counterTwoPixelStream_s2mPipe_ready) begin
      compareStage_counterTwoPixelStream_s2mPipe_rData <= compareStage_counterTwoPixelStream_s2mPipe_payload;
    end
    if(compareStage_mainThreePixelStream_ready) begin
      compareStage_mainThreePixelStream_rData <= compareStage_mainThreePixelStream_payload;
    end
    if(compareStage_mainThreePixelStream_s2mPipe_ready) begin
      compareStage_mainThreePixelStream_s2mPipe_rData <= compareStage_mainThreePixelStream_s2mPipe_payload;
    end
    if(compareStage_counterThreePixelStream_ready) begin
      compareStage_counterThreePixelStream_rData <= compareStage_counterThreePixelStream_payload;
    end
    if(compareStage_counterThreePixelStream_s2mPipe_ready) begin
      compareStage_counterThreePixelStream_s2mPipe_rData <= compareStage_counterThreePixelStream_s2mPipe_payload;
    end
    if(compareStage_mainOneValidStream_ready) begin
      compareStage_mainOneValidStream_rData <= compareStage_mainOneValidStream_payload;
    end
    if(compareStage_mainOneValidStream_s2mPipe_ready) begin
      compareStage_mainOneValidStream_s2mPipe_rData <= compareStage_mainOneValidStream_s2mPipe_payload;
    end
    if(compareStage_counterOneValidStream_ready) begin
      compareStage_counterOneValidStream_rData <= compareStage_counterOneValidStream_payload;
    end
    if(compareStage_counterOneValidStream_s2mPipe_ready) begin
      compareStage_counterOneValidStream_s2mPipe_rData <= compareStage_counterOneValidStream_s2mPipe_payload;
    end
    if(compareStage_mainTwoValidStream_ready) begin
      compareStage_mainTwoValidStream_rData <= compareStage_mainTwoValidStream_payload;
    end
    if(compareStage_mainTwoValidStream_s2mPipe_ready) begin
      compareStage_mainTwoValidStream_s2mPipe_rData <= compareStage_mainTwoValidStream_s2mPipe_payload;
    end
    if(compareStage_counterTwoValidStream_ready) begin
      compareStage_counterTwoValidStream_rData <= compareStage_counterTwoValidStream_payload;
    end
    if(compareStage_counterTwoValidStream_s2mPipe_ready) begin
      compareStage_counterTwoValidStream_s2mPipe_rData <= compareStage_counterTwoValidStream_s2mPipe_payload;
    end
    if(compareStage_mainThreeValidStream_ready) begin
      compareStage_mainThreeValidStream_rData <= compareStage_mainThreeValidStream_payload;
    end
    if(compareStage_mainThreeValidStream_s2mPipe_ready) begin
      compareStage_mainThreeValidStream_s2mPipe_rData <= compareStage_mainThreeValidStream_s2mPipe_payload;
    end
    if(compareStage_counterThreeValidStream_ready) begin
      compareStage_counterThreeValidStream_rData <= compareStage_counterThreeValidStream_payload;
    end
    if(compareStage_counterThreeValidStream_s2mPipe_ready) begin
      compareStage_counterThreeValidStream_s2mPipe_rData <= compareStage_counterThreeValidStream_s2mPipe_payload;
    end
    if(compareStage_controlPipe_translated_ready) begin
      compareStage_controlPipe_translated_rData_frameStart <= compareStage_controlPipe_translated_payload_frameStart;
      compareStage_controlPipe_translated_rData_rowEnd <= compareStage_controlPipe_translated_payload_rowEnd;
      compareStage_controlPipe_translated_rData_pipeValid <= compareStage_controlPipe_translated_payload_pipeValid;
      compareStage_controlPipe_translated_rData_firstRow <= compareStage_controlPipe_translated_payload_firstRow;
      compareStage_controlPipe_translated_rData_lastRow <= compareStage_controlPipe_translated_payload_lastRow;
      compareStage_controlPipe_translated_rData_finalResult <= compareStage_controlPipe_translated_payload_finalResult;
      compareStage_controlPipe_translated_rData_mainCompare <= compareStage_controlPipe_translated_payload_mainCompare;
      compareStage_controlPipe_translated_rData_counterCompare <= compareStage_controlPipe_translated_payload_counterCompare;
      compareStage_controlPipe_translated_rData_horizontalCompare <= compareStage_controlPipe_translated_payload_horizontalCompare;
      compareStage_controlPipe_translated_rData_verticalCompare <= compareStage_controlPipe_translated_payload_verticalCompare;
      compareStage_controlPipe_translated_rData_mainDiff <= compareStage_controlPipe_translated_payload_mainDiff;
      compareStage_controlPipe_translated_rData_counterDiff <= compareStage_controlPipe_translated_payload_counterDiff;
      compareStage_controlPipe_translated_rData_horizontalDiff <= compareStage_controlPipe_translated_payload_horizontalDiff;
      compareStage_controlPipe_translated_rData_verticalDiff <= compareStage_controlPipe_translated_payload_verticalDiff;
      compareStage_controlPipe_translated_rData_isHorizontalMin <= compareStage_controlPipe_translated_payload_isHorizontalMin;
      compareStage_controlPipe_translated_rData_minDiff <= compareStage_controlPipe_translated_payload_minDiff;
      compareStage_controlPipe_translated_rData_currentPosition <= compareStage_controlPipe_translated_payload_currentPosition;
      compareStage_controlPipe_translated_rData_nextPosition <= compareStage_controlPipe_translated_payload_nextPosition;
      compareStage_controlPipe_translated_rData_horizontalDirectionValid <= compareStage_controlPipe_translated_payload_horizontalDirectionValid;
      compareStage_controlPipe_translated_rData_verticalDirectionValid <= compareStage_controlPipe_translated_payload_verticalDirectionValid;
      compareStage_controlPipe_translated_rData_mainDirectionValid <= compareStage_controlPipe_translated_payload_mainDirectionValid;
      compareStage_controlPipe_translated_rData_counterDirectionValid <= compareStage_controlPipe_translated_payload_counterDirectionValid;
      compareStage_controlPipe_translated_rData_inValidMinDiff <= compareStage_controlPipe_translated_payload_inValidMinDiff;
    end
    if(compareStage_controlPipe_translated_s2mPipe_ready) begin
      compareStage_controlPipe_translated_s2mPipe_rData_frameStart <= compareStage_controlPipe_translated_s2mPipe_payload_frameStart;
      compareStage_controlPipe_translated_s2mPipe_rData_rowEnd <= compareStage_controlPipe_translated_s2mPipe_payload_rowEnd;
      compareStage_controlPipe_translated_s2mPipe_rData_pipeValid <= compareStage_controlPipe_translated_s2mPipe_payload_pipeValid;
      compareStage_controlPipe_translated_s2mPipe_rData_firstRow <= compareStage_controlPipe_translated_s2mPipe_payload_firstRow;
      compareStage_controlPipe_translated_s2mPipe_rData_lastRow <= compareStage_controlPipe_translated_s2mPipe_payload_lastRow;
      compareStage_controlPipe_translated_s2mPipe_rData_finalResult <= compareStage_controlPipe_translated_s2mPipe_payload_finalResult;
      compareStage_controlPipe_translated_s2mPipe_rData_mainCompare <= compareStage_controlPipe_translated_s2mPipe_payload_mainCompare;
      compareStage_controlPipe_translated_s2mPipe_rData_counterCompare <= compareStage_controlPipe_translated_s2mPipe_payload_counterCompare;
      compareStage_controlPipe_translated_s2mPipe_rData_horizontalCompare <= compareStage_controlPipe_translated_s2mPipe_payload_horizontalCompare;
      compareStage_controlPipe_translated_s2mPipe_rData_verticalCompare <= compareStage_controlPipe_translated_s2mPipe_payload_verticalCompare;
      compareStage_controlPipe_translated_s2mPipe_rData_mainDiff <= compareStage_controlPipe_translated_s2mPipe_payload_mainDiff;
      compareStage_controlPipe_translated_s2mPipe_rData_counterDiff <= compareStage_controlPipe_translated_s2mPipe_payload_counterDiff;
      compareStage_controlPipe_translated_s2mPipe_rData_horizontalDiff <= compareStage_controlPipe_translated_s2mPipe_payload_horizontalDiff;
      compareStage_controlPipe_translated_s2mPipe_rData_verticalDiff <= compareStage_controlPipe_translated_s2mPipe_payload_verticalDiff;
      compareStage_controlPipe_translated_s2mPipe_rData_isHorizontalMin <= compareStage_controlPipe_translated_s2mPipe_payload_isHorizontalMin;
      compareStage_controlPipe_translated_s2mPipe_rData_minDiff <= compareStage_controlPipe_translated_s2mPipe_payload_minDiff;
      compareStage_controlPipe_translated_s2mPipe_rData_currentPosition <= compareStage_controlPipe_translated_s2mPipe_payload_currentPosition;
      compareStage_controlPipe_translated_s2mPipe_rData_nextPosition <= compareStage_controlPipe_translated_s2mPipe_payload_nextPosition;
      compareStage_controlPipe_translated_s2mPipe_rData_horizontalDirectionValid <= compareStage_controlPipe_translated_s2mPipe_payload_horizontalDirectionValid;
      compareStage_controlPipe_translated_s2mPipe_rData_verticalDirectionValid <= compareStage_controlPipe_translated_s2mPipe_payload_verticalDirectionValid;
      compareStage_controlPipe_translated_s2mPipe_rData_mainDirectionValid <= compareStage_controlPipe_translated_s2mPipe_payload_mainDirectionValid;
      compareStage_controlPipe_translated_s2mPipe_rData_counterDirectionValid <= compareStage_controlPipe_translated_s2mPipe_payload_counterDirectionValid;
      compareStage_controlPipe_translated_s2mPipe_rData_inValidMinDiff <= compareStage_controlPipe_translated_s2mPipe_payload_inValidMinDiff;
    end
    if(diffStage_mainOnePixelStream_ready) begin
      diffStage_mainOnePixelStream_rData <= diffStage_mainOnePixelStream_payload;
    end
    if(diffStage_mainOnePixelStream_s2mPipe_ready) begin
      diffStage_mainOnePixelStream_s2mPipe_rData <= diffStage_mainOnePixelStream_s2mPipe_payload;
    end
    if(diffStage_counterOnePixelStream_ready) begin
      diffStage_counterOnePixelStream_rData <= diffStage_counterOnePixelStream_payload;
    end
    if(diffStage_counterOnePixelStream_s2mPipe_ready) begin
      diffStage_counterOnePixelStream_s2mPipe_rData <= diffStage_counterOnePixelStream_s2mPipe_payload;
    end
    if(diffStage_mainTwoPixelStream_ready) begin
      diffStage_mainTwoPixelStream_rData <= diffStage_mainTwoPixelStream_payload;
    end
    if(diffStage_mainTwoPixelStream_s2mPipe_ready) begin
      diffStage_mainTwoPixelStream_s2mPipe_rData <= diffStage_mainTwoPixelStream_s2mPipe_payload;
    end
    if(diffStage_counterTwoPixelStream_ready) begin
      diffStage_counterTwoPixelStream_rData <= diffStage_counterTwoPixelStream_payload;
    end
    if(diffStage_counterTwoPixelStream_s2mPipe_ready) begin
      diffStage_counterTwoPixelStream_s2mPipe_rData <= diffStage_counterTwoPixelStream_s2mPipe_payload;
    end
    if(diffStage_mainThreePixelStream_ready) begin
      diffStage_mainThreePixelStream_rData <= diffStage_mainThreePixelStream_payload;
    end
    if(diffStage_mainThreePixelStream_s2mPipe_ready) begin
      diffStage_mainThreePixelStream_s2mPipe_rData <= diffStage_mainThreePixelStream_s2mPipe_payload;
    end
    if(diffStage_counterThreePixelStream_ready) begin
      diffStage_counterThreePixelStream_rData <= diffStage_counterThreePixelStream_payload;
    end
    if(diffStage_counterThreePixelStream_s2mPipe_ready) begin
      diffStage_counterThreePixelStream_s2mPipe_rData <= diffStage_counterThreePixelStream_s2mPipe_payload;
    end
    if(diffStage_mainOneValidStream_ready) begin
      diffStage_mainOneValidStream_rData <= diffStage_mainOneValidStream_payload;
    end
    if(diffStage_mainOneValidStream_s2mPipe_ready) begin
      diffStage_mainOneValidStream_s2mPipe_rData <= diffStage_mainOneValidStream_s2mPipe_payload;
    end
    if(diffStage_counterOneValidStream_ready) begin
      diffStage_counterOneValidStream_rData <= diffStage_counterOneValidStream_payload;
    end
    if(diffStage_counterOneValidStream_s2mPipe_ready) begin
      diffStage_counterOneValidStream_s2mPipe_rData <= diffStage_counterOneValidStream_s2mPipe_payload;
    end
    if(diffStage_mainTwoValidStream_ready) begin
      diffStage_mainTwoValidStream_rData <= diffStage_mainTwoValidStream_payload;
    end
    if(diffStage_mainTwoValidStream_s2mPipe_ready) begin
      diffStage_mainTwoValidStream_s2mPipe_rData <= diffStage_mainTwoValidStream_s2mPipe_payload;
    end
    if(diffStage_counterTwoValidStream_ready) begin
      diffStage_counterTwoValidStream_rData <= diffStage_counterTwoValidStream_payload;
    end
    if(diffStage_counterTwoValidStream_s2mPipe_ready) begin
      diffStage_counterTwoValidStream_s2mPipe_rData <= diffStage_counterTwoValidStream_s2mPipe_payload;
    end
    if(diffStage_mainThreeValidStream_ready) begin
      diffStage_mainThreeValidStream_rData <= diffStage_mainThreeValidStream_payload;
    end
    if(diffStage_mainThreeValidStream_s2mPipe_ready) begin
      diffStage_mainThreeValidStream_s2mPipe_rData <= diffStage_mainThreeValidStream_s2mPipe_payload;
    end
    if(diffStage_counterThreeValidStream_ready) begin
      diffStage_counterThreeValidStream_rData <= diffStage_counterThreeValidStream_payload;
    end
    if(diffStage_counterThreeValidStream_s2mPipe_ready) begin
      diffStage_counterThreeValidStream_s2mPipe_rData <= diffStage_counterThreeValidStream_s2mPipe_payload;
    end
    if(resultStage_controlPipeBeforePipe_ready) begin
      resultStage_controlPipeBeforePipe_rData_frameStart <= resultStage_controlPipeBeforePipe_payload_frameStart;
      resultStage_controlPipeBeforePipe_rData_rowEnd <= resultStage_controlPipeBeforePipe_payload_rowEnd;
      resultStage_controlPipeBeforePipe_rData_pipeValid <= resultStage_controlPipeBeforePipe_payload_pipeValid;
      resultStage_controlPipeBeforePipe_rData_firstRow <= resultStage_controlPipeBeforePipe_payload_firstRow;
      resultStage_controlPipeBeforePipe_rData_lastRow <= resultStage_controlPipeBeforePipe_payload_lastRow;
      resultStage_controlPipeBeforePipe_rData_finalResult <= resultStage_controlPipeBeforePipe_payload_finalResult;
      resultStage_controlPipeBeforePipe_rData_mainCompare <= resultStage_controlPipeBeforePipe_payload_mainCompare;
      resultStage_controlPipeBeforePipe_rData_counterCompare <= resultStage_controlPipeBeforePipe_payload_counterCompare;
      resultStage_controlPipeBeforePipe_rData_horizontalCompare <= resultStage_controlPipeBeforePipe_payload_horizontalCompare;
      resultStage_controlPipeBeforePipe_rData_verticalCompare <= resultStage_controlPipeBeforePipe_payload_verticalCompare;
      resultStage_controlPipeBeforePipe_rData_mainDiff <= resultStage_controlPipeBeforePipe_payload_mainDiff;
      resultStage_controlPipeBeforePipe_rData_counterDiff <= resultStage_controlPipeBeforePipe_payload_counterDiff;
      resultStage_controlPipeBeforePipe_rData_horizontalDiff <= resultStage_controlPipeBeforePipe_payload_horizontalDiff;
      resultStage_controlPipeBeforePipe_rData_verticalDiff <= resultStage_controlPipeBeforePipe_payload_verticalDiff;
      resultStage_controlPipeBeforePipe_rData_isHorizontalMin <= resultStage_controlPipeBeforePipe_payload_isHorizontalMin;
      resultStage_controlPipeBeforePipe_rData_minDiff <= resultStage_controlPipeBeforePipe_payload_minDiff;
      resultStage_controlPipeBeforePipe_rData_currentPosition <= resultStage_controlPipeBeforePipe_payload_currentPosition;
      resultStage_controlPipeBeforePipe_rData_nextPosition <= resultStage_controlPipeBeforePipe_payload_nextPosition;
      resultStage_controlPipeBeforePipe_rData_horizontalDirectionValid <= resultStage_controlPipeBeforePipe_payload_horizontalDirectionValid;
      resultStage_controlPipeBeforePipe_rData_verticalDirectionValid <= resultStage_controlPipeBeforePipe_payload_verticalDirectionValid;
      resultStage_controlPipeBeforePipe_rData_mainDirectionValid <= resultStage_controlPipeBeforePipe_payload_mainDirectionValid;
      resultStage_controlPipeBeforePipe_rData_counterDirectionValid <= resultStage_controlPipeBeforePipe_payload_counterDirectionValid;
      resultStage_controlPipeBeforePipe_rData_inValidMinDiff <= resultStage_controlPipeBeforePipe_payload_inValidMinDiff;
    end
    if(resultStage_controlPipeBeforePipe_s2mPipe_ready) begin
      resultStage_controlPipeBeforePipe_s2mPipe_rData_frameStart <= resultStage_controlPipeBeforePipe_s2mPipe_payload_frameStart;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_rowEnd <= resultStage_controlPipeBeforePipe_s2mPipe_payload_rowEnd;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_pipeValid <= resultStage_controlPipeBeforePipe_s2mPipe_payload_pipeValid;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_firstRow <= resultStage_controlPipeBeforePipe_s2mPipe_payload_firstRow;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_lastRow <= resultStage_controlPipeBeforePipe_s2mPipe_payload_lastRow;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_finalResult <= resultStage_controlPipeBeforePipe_s2mPipe_payload_finalResult;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_mainCompare <= resultStage_controlPipeBeforePipe_s2mPipe_payload_mainCompare;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_counterCompare <= resultStage_controlPipeBeforePipe_s2mPipe_payload_counterCompare;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_horizontalCompare <= resultStage_controlPipeBeforePipe_s2mPipe_payload_horizontalCompare;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_verticalCompare <= resultStage_controlPipeBeforePipe_s2mPipe_payload_verticalCompare;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_mainDiff <= resultStage_controlPipeBeforePipe_s2mPipe_payload_mainDiff;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_counterDiff <= resultStage_controlPipeBeforePipe_s2mPipe_payload_counterDiff;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_horizontalDiff <= resultStage_controlPipeBeforePipe_s2mPipe_payload_horizontalDiff;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_verticalDiff <= resultStage_controlPipeBeforePipe_s2mPipe_payload_verticalDiff;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_isHorizontalMin <= resultStage_controlPipeBeforePipe_s2mPipe_payload_isHorizontalMin;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_minDiff <= resultStage_controlPipeBeforePipe_s2mPipe_payload_minDiff;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_currentPosition <= resultStage_controlPipeBeforePipe_s2mPipe_payload_currentPosition;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_nextPosition <= resultStage_controlPipeBeforePipe_s2mPipe_payload_nextPosition;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_horizontalDirectionValid <= resultStage_controlPipeBeforePipe_s2mPipe_payload_horizontalDirectionValid;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_verticalDirectionValid <= resultStage_controlPipeBeforePipe_s2mPipe_payload_verticalDirectionValid;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_mainDirectionValid <= resultStage_controlPipeBeforePipe_s2mPipe_payload_mainDirectionValid;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_counterDirectionValid <= resultStage_controlPipeBeforePipe_s2mPipe_payload_counterDirectionValid;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_inValidMinDiff <= resultStage_controlPipeBeforePipe_s2mPipe_payload_inValidMinDiff;
    end
    if(resultStage_pixelStream_ready) begin
      resultStage_pixelStream_rData <= resultStage_pixelStream_payload;
    end
    if(resultStage_pixelStream_s2mPipe_ready) begin
      resultStage_pixelStream_s2mPipe_rData <= resultStage_pixelStream_s2mPipe_payload;
    end
    if(pixelsStream_ready) begin
      pixelsStream_rData_pixel <= pixelsStream_payload_pixel;
      pixelsStream_rData_frameStart <= pixelsStream_payload_frameStart;
      pixelsStream_rData_rowEnd <= pixelsStream_payload_rowEnd;
    end
    if(pixelsStream_s2mPipe_ready) begin
      pixelsStream_s2mPipe_rData_pixel <= pixelsStream_s2mPipe_payload_pixel;
      pixelsStream_s2mPipe_rData_frameStart <= pixelsStream_s2mPipe_payload_frameStart;
      pixelsStream_s2mPipe_rData_rowEnd <= pixelsStream_s2mPipe_payload_rowEnd;
    end
  end


endmodule

module SuperResolutionPart2_2 (
  input               pixelsIn_valid,
  output reg          pixelsIn_ready,
  input      [7:0]    pixelsIn_payload_pixel,
  input               pixelsIn_payload_frameStart,
  input               pixelsIn_payload_rowEnd,
  input               startIn,
  input               inpThreeDoneIn,
  output reg          pixelsOut_valid,
  input               pixelsOut_ready,
  output reg [7:0]    pixelsOut_payload_pixel,
  output reg          pixelsOut_payload_frameStart,
  output reg          pixelsOut_payload_rowEnd,
  output reg          pixelsOut_payload_inpValid,
  output reg          startOut,
  output reg          inpTwoDoneOut,
  input      [7:0]    thresholdIn,
  input      [9:0]    widthIn,
  input      [9:0]    heightIn,
  input               clk,
  input               resetn
);
  localparam controlStateMachine_enumDef_7_BOOT = 3'd0;
  localparam controlStateMachine_enumDef_7_HOLD = 3'd1;
  localparam controlStateMachine_enumDef_7_PASS = 3'd2;
  localparam controlStateMachine_enumDef_7_ONCE = 3'd3;
  localparam controlStateMachine_enumDef_7_TWICE = 3'd4;

  reg        [7:0]    CICC1851_lineBufferOne_port1;
  reg        [7:0]    CICC1851_lineBufferOne_port2;
  reg        [7:0]    CICC1851_lineBufferTwo_port1;
  reg        [7:0]    CICC1851_lineBufferTwo_port2;
  reg        [7:0]    CICC1851_lineBufferOdd_port1;
  wire                diffStage_controlPipe_fork_io_input_ready;
  wire                diffStage_controlPipe_fork_io_outputs_0_valid;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_frameStart;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_rowEnd;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_passMode;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_passValid;
  wire       [2:0]    diffStage_controlPipe_fork_io_outputs_0_payload_onceMode;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_onceValid;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_mainCompare;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_counterCompare;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_payload_mainDiff;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_payload_counterDiff;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_twiceCompValid;
  wire       [2:0]    diffStage_controlPipe_fork_io_outputs_0_payload_twiceMode;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_inpValidFlag;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_oddValid;
  wire                diffStage_controlPipe_fork_io_outputs_1_valid;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_frameStart;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_rowEnd;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_passMode;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_passValid;
  wire       [2:0]    diffStage_controlPipe_fork_io_outputs_1_payload_onceMode;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_onceValid;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_mainCompare;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_counterCompare;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_twiceCompValid;
  wire       [2:0]    diffStage_controlPipe_fork_io_outputs_1_payload_twiceMode;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_inpValidFlag;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_oddValid;
  wire       [10:0]   CICC1851_bufferRowCount_valueNext;
  wire       [0:0]    CICC1851_bufferRowCount_valueNext_1;
  wire       [10:0]   CICC1851_bufferWAddr_valueNext;
  wire       [0:0]    CICC1851_bufferWAddr_valueNext_1;
  wire       [11:0]   CICC1851_outPixelAddr_valueNext;
  wire       [0:0]    CICC1851_outPixelAddr_valueNext_1;
  wire       [11:0]   CICC1851_outRowCount_valueNext;
  wire       [0:0]    CICC1851_outRowCount_valueNext_1;
  wire       [11:0]   CICC1851_alreadySendRow_valueNext;
  wire       [0:0]    CICC1851_alreadySendRow_valueNext_1;
  wire       [11:0]   CICC1851_alreadySendCountInRow_valueNext;
  wire       [0:0]    CICC1851_alreadySendCountInRow_valueNext_1;
  wire       [11:0]   CICC1851_mainAddrOne;
  wire       [11:0]   CICC1851_counterAddrOne;
  wire       [11:0]   CICC1851_mainAddrTwo;
  wire       [11:0]   CICC1851_counterAddrTwo;
  wire       [11:0]   CICC1851_oddAddr;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l181;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l181_1;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l181_2;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l182;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l182_1;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l182_2;
  wire       [10:0]   CICC1851_when_SuperResolutionPart2_l195;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l218;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l234;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l234_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l234_2;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l235;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l235_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l235_2;
  wire       [7:0]    CICC1851_lineBufferOne_port;
  wire                CICC1851_lineBufferOne_port_1;
  wire       [7:0]    CICC1851_lineBufferOdd_port;
  wire                CICC1851_lineBufferOdd_port_1;
  wire       [7:0]    CICC1851_lineBufferTwo_port;
  wire                CICC1851_lineBufferTwo_port_1;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_1;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_2;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_3;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_4;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_5;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_6;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_7;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_8;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_9;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_10;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_11;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_12;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_13;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_14;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_15;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_16;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_17;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_18;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_19;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l763;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l763_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l763_2;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l764;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l764_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l764_2;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l783;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l785;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l787;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l789;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l793;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l796;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l799;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l802;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l560;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l560_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l602;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l602_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l602_2;
  wire       [2:0]    CICC1851_when_SuperResolutionPart2_l602_3;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l603;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l603_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l605;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l605_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l605_2;
  wire       [2:0]    CICC1851_when_SuperResolutionPart2_l605_3;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l606;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l606_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l606_2;
  wire       [1:0]    CICC1851_when_SuperResolutionPart2_l606_3;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l609;
  wire       [11:0]   CICC1851_mainAddrOne_1;
  wire       [11:0]   CICC1851_mainAddrOne_2;
  wire       [11:0]   CICC1851_mainAddrTwo_1;
  wire       [11:0]   CICC1851_mainAddrTwo_2;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l667;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l667_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l667_2;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l667_3;
  wire       [1:0]    CICC1851_when_SuperResolutionPart2_l667_4;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l668;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l668_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l668_2;
  wire       [1:0]    CICC1851_when_SuperResolutionPart2_l668_3;
  wire       [11:0]   CICC1851_mainAddrOne_3;
  wire       [11:0]   CICC1851_mainAddrOne_4;
  wire       [11:0]   CICC1851_mainAddrTwo_3;
  wire       [11:0]   CICC1851_mainAddrTwo_4;
  wire       [1:0]    CICC1851_controls_onceMode;
  wire       [1:0]    CICC1851_controls_onceMode_1;
  wire       [11:0]   CICC1851_mainAddrOne_5;
  wire       [11:0]   CICC1851_mainAddrOne_6;
  wire       [11:0]   CICC1851_counterAddrOne_1;
  wire       [11:0]   CICC1851_counterAddrOne_2;
  wire       [11:0]   CICC1851_counterAddrOne_3;
  wire       [11:0]   CICC1851_counterAddrOne_4;
  wire       [0:0]    CICC1851_controls_onceMode_2;
  wire       [11:0]   CICC1851_mainAddrTwo_5;
  wire       [11:0]   CICC1851_mainAddrTwo_6;
  wire       [11:0]   CICC1851_counterAddrTwo_1;
  wire       [11:0]   CICC1851_counterAddrTwo_2;
  wire       [11:0]   CICC1851_counterAddrTwo_3;
  wire       [11:0]   CICC1851_counterAddrTwo_4;
  wire       [11:0]   CICC1851_mainAddrOne_7;
  wire       [11:0]   CICC1851_mainAddrOne_8;
  wire       [11:0]   CICC1851_mainAddrOne_9;
  wire       [11:0]   CICC1851_mainAddrOne_10;
  wire       [12:0]   CICC1851_counterAddrOne_5;
  wire       [12:0]   CICC1851_counterAddrOne_6;
  wire       [12:0]   CICC1851_counterAddrOne_7;
  wire       [1:0]    CICC1851_counterAddrOne_8;
  wire       [1:0]    CICC1851_controls_twiceMode;
  wire       [11:0]   CICC1851_mainAddrTwo_7;
  wire       [11:0]   CICC1851_mainAddrTwo_8;
  wire       [1:0]    CICC1851_controls_twiceMode_1;
  wire       [11:0]   CICC1851_mainAddrTwo_9;
  wire       [11:0]   CICC1851_mainAddrTwo_10;
  wire       [12:0]   CICC1851_counterAddrTwo_5;
  wire       [12:0]   CICC1851_counterAddrTwo_6;
  wire       [12:0]   CICC1851_counterAddrTwo_7;
  wire       [1:0]    CICC1851_counterAddrTwo_8;
  wire       [11:0]   CICC1851_mainAddrOne_11;
  wire       [11:0]   CICC1851_mainAddrOne_12;
  wire       [11:0]   CICC1851_counterAddrTwo_9;
  wire       [11:0]   CICC1851_counterAddrTwo_10;
  wire       [11:0]   CICC1851_mainAddrTwo_11;
  wire       [11:0]   CICC1851_mainAddrTwo_12;
  wire       [11:0]   CICC1851_counterAddrOne_9;
  wire       [11:0]   CICC1851_counterAddrOne_10;
  wire       [12:0]   CICC1851_mainAddrTwo_13;
  wire       [12:0]   CICC1851_mainAddrTwo_14;
  wire       [12:0]   CICC1851_mainAddrTwo_15;
  wire       [1:0]    CICC1851_mainAddrTwo_16;
  wire       [12:0]   CICC1851_counterAddrOne_11;
  wire       [12:0]   CICC1851_counterAddrOne_12;
  wire       [12:0]   CICC1851_counterAddrOne_13;
  wire       [1:0]    CICC1851_counterAddrOne_14;
  wire       [0:0]    CICC1851_controls_twiceMode_2;
  wire       [11:0]   CICC1851_mainAddrTwo_17;
  wire       [11:0]   CICC1851_mainAddrTwo_18;
  wire       [11:0]   CICC1851_counterAddrOne_15;
  wire       [11:0]   CICC1851_counterAddrOne_16;
  wire       [11:0]   CICC1851_mainAddrOne_13;
  wire       [11:0]   CICC1851_mainAddrOne_14;
  wire       [11:0]   CICC1851_counterAddrTwo_11;
  wire       [11:0]   CICC1851_counterAddrTwo_12;
  wire       [12:0]   CICC1851_mainAddrOne_15;
  wire       [12:0]   CICC1851_mainAddrOne_16;
  wire       [12:0]   CICC1851_mainAddrOne_17;
  wire       [1:0]    CICC1851_mainAddrOne_18;
  wire       [12:0]   CICC1851_counterAddrTwo_13;
  wire       [12:0]   CICC1851_counterAddrTwo_14;
  wire       [12:0]   CICC1851_counterAddrTwo_15;
  wire       [1:0]    CICC1851_counterAddrTwo_16;
  reg                 inpTwoDone;
  reg                 startIn_regNext;
  wire                when_SuperResolutionPart2_l40;
  reg                 readDone;
  wire                when_SuperResolutionPart2_l43;
  reg                 startRead;
  wire                when_SuperResolutionPart2_l46;
  wire                when_SuperResolutionPart2_l46_1;
  reg                 slaveStart;
  wire                pixelsIn_fire;
  wire                when_SuperResolutionPart2_l49;
  wire                when_SuperResolutionPart2_l49_1;
  reg                 frameStart;
  reg        [7:0]    inpThreshold;
  reg        [9:0]    bmpWidth;
  reg        [9:0]    bmpHeight;
  reg                 holdBuffer;
  wire                when_SuperResolutionPart2_l64;
  reg                 writeDone;
  wire                when_SuperResolutionPart2_l67;
  reg                 bufferRowCount_willIncrement;
  reg                 bufferRowCount_willClear;
  reg        [10:0]   bufferRowCount_valueNext;
  reg        [10:0]   bufferRowCount_value;
  wire                bufferRowCount_willOverflowIfInc;
  wire                bufferRowCount_willOverflow;
  reg                 bufferReuse;
  reg                 bufferEnable;
  wire                when_SuperResolutionPart2_l76;
  wire                when_SuperResolutionPart2_l76_1;
  reg        [1:0]    bufferSwitch;
  reg                 nextRowBuffer;
  wire                when_SuperResolutionPart2_l82;
  reg                 bufferWAddr_willIncrement;
  reg                 bufferWAddr_willClear;
  reg        [10:0]   bufferWAddr_valueNext;
  reg        [10:0]   bufferWAddr_value;
  wire                bufferWAddr_willOverflowIfInc;
  wire                bufferWAddr_willOverflow;
  reg                 outPixelAddr_willIncrement;
  reg                 outPixelAddr_willClear;
  reg        [11:0]   outPixelAddr_valueNext;
  reg        [11:0]   outPixelAddr_value;
  wire                outPixelAddr_willOverflowIfInc;
  wire                outPixelAddr_willOverflow;
  reg                 outRowCount_willIncrement;
  reg                 outRowCount_willClear;
  reg        [11:0]   outRowCount_valueNext;
  reg        [11:0]   outRowCount_value;
  wire                outRowCount_willOverflowIfInc;
  wire                outRowCount_willOverflow;
  reg                 alreadySendRow_willIncrement;
  reg                 alreadySendRow_willClear;
  reg        [11:0]   alreadySendRow_valueNext;
  reg        [11:0]   alreadySendRow_value;
  wire                alreadySendRow_willOverflowIfInc;
  wire                alreadySendRow_willOverflow;
  reg                 alreadySendCountInRow_willIncrement;
  reg                 alreadySendCountInRow_willClear;
  reg        [11:0]   alreadySendCountInRow_valueNext;
  reg        [11:0]   alreadySendCountInRow_value;
  wire                alreadySendCountInRow_willOverflowIfInc;
  wire                alreadySendCountInRow_willOverflow;
  reg                 alreadyReachRowEnd;
  reg                 alreadyReachFinalRow;
  reg                 outReachRowEnd;
  reg                 outReachFinalRow;
  reg                 bufferReachRowEnd;
  reg                 bufferReachFinalRow;
  reg                 oddBufferRow;
  reg                 startIn_regNext_1;
  wire                when_SuperResolutionPart2_l106;
  reg                 zeroInFourOutPixelAddr;
  reg                 startIn_regNext_2;
  wire                when_SuperResolutionPart2_l108;
  reg                 oneInFourOutPixelAddr;
  reg                 startIn_regNext_3;
  wire                when_SuperResolutionPart2_l109;
  reg                 twoInFourOutPixelAddr;
  reg                 startIn_regNext_4;
  wire                when_SuperResolutionPart2_l110;
  reg                 threeInFourOutPixelAddr;
  reg                 startIn_regNext_5;
  wire                when_SuperResolutionPart2_l111;
  reg                 zeroInFourOutRow;
  reg                 startIn_regNext_6;
  wire                when_SuperResolutionPart2_l113;
  reg                 oneInFourOutRow;
  reg                 startIn_regNext_7;
  wire                when_SuperResolutionPart2_l114;
  reg                 twoInFourOutRow;
  reg                 startIn_regNext_8;
  wire                when_SuperResolutionPart2_l115;
  reg                 threeInFourOutRow;
  reg                 startIn_regNext_9;
  wire                when_SuperResolutionPart2_l116;
  wire       [2:0]    currentState;
  reg                 willHoldToTwice;
  reg                 startIn_regNext_10;
  wire                when_SuperResolutionPart2_l120;
  reg                 willPassToHoldCaseOne;
  reg                 startIn_regNext_11;
  wire                when_SuperResolutionPart2_l121;
  reg                 willPassToHoldCaseTwo;
  reg                 startIn_regNext_12;
  wire                when_SuperResolutionPart2_l122;
  reg                 holdWillPassToHoldCaseTwo;
  reg                 startIn_regNext_13;
  wire                when_SuperResolutionPart2_l123;
  reg                 willOnceToHoldCaseOne;
  reg                 startIn_regNext_14;
  wire                when_SuperResolutionPart2_l124;
  reg                 willOnceToHoldCaseTwo;
  reg                 startIn_regNext_15;
  wire                when_SuperResolutionPart2_l125;
  reg                 willOnceToHoldCaseThree;
  reg                 startIn_regNext_16;
  wire                when_SuperResolutionPart2_l126;
  wire                when_SuperResolutionPart2_l134;
  reg        [10:0]   mainAddrOne;
  reg        [10:0]   counterAddrOne;
  reg        [10:0]   mainAddrTwo;
  reg        [10:0]   counterAddrTwo;
  wire       [10:0]   oddAddr;
  wire                validStream_valid;
  reg                 validStream_ready;
  wire                controlStream_valid;
  wire                controlStream_ready;
  wire                controlStream_payload_frameStart;
  wire                controlStream_payload_rowEnd;
  wire                controlStream_payload_passMode;
  wire                controlStream_payload_passValid;
  wire       [2:0]    controlStream_payload_onceMode;
  wire                controlStream_payload_onceValid;
  wire                controlStream_payload_mainCompare;
  wire                controlStream_payload_counterCompare;
  wire       [7:0]    controlStream_payload_mainDiff;
  wire       [7:0]    controlStream_payload_counterDiff;
  wire                controlStream_payload_twiceCompValid;
  wire       [2:0]    controlStream_payload_twiceMode;
  wire                controlStream_payload_inpValidFlag;
  wire                controlStream_payload_oddValid;
  reg                 controls_frameStart;
  reg                 controls_rowEnd;
  reg                 controls_passMode;
  reg                 controls_passValid;
  reg        [2:0]    controls_onceMode;
  reg                 controls_onceValid;
  wire                controls_mainCompare;
  wire                controls_counterCompare;
  wire       [7:0]    controls_mainDiff;
  wire       [7:0]    controls_counterDiff;
  reg                 controls_twiceCompValid;
  reg        [2:0]    controls_twiceMode;
  reg                 controls_inpValidFlag;
  reg                 controls_oddValid;
  wire       [31:0]   CICC1851_controls_frameStart;
  wire                mainAddrOneStream_valid;
  wire                mainAddrOneStream_ready;
  wire       [10:0]   mainAddrOneStream_payload;
  wire                counterAddrOneStream_valid;
  wire                counterAddrOneStream_ready;
  wire       [10:0]   counterAddrOneStream_payload;
  wire                mainAddrTwoStream_valid;
  wire                mainAddrTwoStream_ready;
  wire       [10:0]   mainAddrTwoStream_payload;
  wire                counterAddrTwoStream_valid;
  wire                counterAddrTwoStream_ready;
  wire       [10:0]   counterAddrTwoStream_payload;
  wire                oddAddrStream_valid;
  wire                oddAddrStream_ready;
  wire       [10:0]   oddAddrStream_payload;
  wire                pixelsIn_s2mPipe_valid;
  reg                 pixelsIn_s2mPipe_ready;
  wire       [7:0]    pixelsIn_s2mPipe_payload_pixel;
  wire                pixelsIn_s2mPipe_payload_frameStart;
  wire                pixelsIn_s2mPipe_payload_rowEnd;
  reg                 pixelsIn_rValid;
  reg        [7:0]    pixelsIn_rData_pixel;
  reg                 pixelsIn_rData_frameStart;
  reg                 pixelsIn_rData_rowEnd;
  wire                pixelsIn_s2mPipe_m2sPipe_valid;
  wire                pixelsIn_s2mPipe_m2sPipe_ready;
  wire       [7:0]    pixelsIn_s2mPipe_m2sPipe_payload_pixel;
  wire                pixelsIn_s2mPipe_m2sPipe_payload_frameStart;
  wire                pixelsIn_s2mPipe_m2sPipe_payload_rowEnd;
  reg                 pixelsIn_s2mPipe_rValid;
  reg        [7:0]    pixelsIn_s2mPipe_rData_pixel;
  reg                 pixelsIn_s2mPipe_rData_frameStart;
  reg                 pixelsIn_s2mPipe_rData_rowEnd;
  wire                when_Stream_l368;
  wire                passPixels_valid;
  wire                passPixels_ready;
  wire       [7:0]    passPixels_payload_pixel;
  wire                passPixels_payload_frameStart;
  wire                passPixels_payload_rowEnd;
  wire                passPixels_fire;
  wire                when_SuperResolutionPart2_l181;
  wire                passPixels_fire_1;
  wire                when_SuperResolutionPart2_l182;
  wire                passPixels_fire_2;
  wire                when_SuperResolutionPart2_l185;
  wire                when_SuperResolutionPart2_l195;
  wire                passPixels_fire_3;
  wire                when_SuperResolutionPart2_l200;
  wire                when_SuperResolutionPart2_l201;
  wire                passPixels_fire_4;
  wire                when_SuperResolutionPart2_l207;
  wire                when_SuperResolutionPart2_l208;
  wire                when_SuperResolutionPart2_l212;
  wire                controlStream_fire;
  wire                when_SuperResolutionPart2_l218;
  wire                when_SuperResolutionPart2_l220;
  wire                passPixels_fire_5;
  wire                when_SuperResolutionPart2_l224;
  wire                pixelsOut_fire;
  wire                when_SuperResolutionPart2_l234;
  wire                pixelsOut_fire_1;
  wire                when_SuperResolutionPart2_l235;
  wire                pixelsOut_fire_2;
  wire                pixelsOut_fire_3;
  wire                when_SuperResolutionPart2_l246;
  wire                passPixels_fire_6;
  wire                passPixels_fire_7;
  wire                passPixels_fire_8;
  wire                passPixels_fire_9;
  wire                passPixels_fire_10;
  wire                controlStream_fire_1;
  wire                pushing;
  wire                passPixels_fire_11;
  wire                controlStream_fire_2;
  wire                poping;
  wire                passPixels_fire_12;
  wire                controlStream_fire_3;
  wire                pushAndPoping;
  wire                mainAddrOneStream_s2mPipe_valid;
  reg                 mainAddrOneStream_s2mPipe_ready;
  wire       [10:0]   mainAddrOneStream_s2mPipe_payload;
  reg                 mainAddrOneStream_rValid;
  reg        [10:0]   mainAddrOneStream_rData;
  wire                mainAddrOneStream_s2mPipe_m2sPipe_valid;
  wire                mainAddrOneStream_s2mPipe_m2sPipe_ready;
  wire       [10:0]   mainAddrOneStream_s2mPipe_m2sPipe_payload;
  reg                 mainAddrOneStream_s2mPipe_rValid;
  reg        [10:0]   mainAddrOneStream_s2mPipe_rData;
  wire                when_Stream_l368_1;
  wire                CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_mainOnePixelStream_payload;
  reg                 CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_1;
  reg                 CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_mainOnePixelStream_payload_1;
  wire                readStage_mainOnePixelStream_valid;
  wire                readStage_mainOnePixelStream_ready;
  wire       [7:0]    readStage_mainOnePixelStream_payload;
  reg                 CICC1851_readStage_mainOnePixelStream_valid;
  reg        [7:0]    CICC1851_readStage_mainOnePixelStream_payload_2;
  wire                when_Stream_l368_2;
  wire                counterAddrOneStream_s2mPipe_valid;
  reg                 counterAddrOneStream_s2mPipe_ready;
  wire       [10:0]   counterAddrOneStream_s2mPipe_payload;
  reg                 counterAddrOneStream_rValid;
  reg        [10:0]   counterAddrOneStream_rData;
  wire                counterAddrOneStream_s2mPipe_m2sPipe_valid;
  wire                counterAddrOneStream_s2mPipe_m2sPipe_ready;
  wire       [10:0]   counterAddrOneStream_s2mPipe_m2sPipe_payload;
  reg                 counterAddrOneStream_s2mPipe_rValid;
  reg        [10:0]   counterAddrOneStream_s2mPipe_rData;
  wire                when_Stream_l368_3;
  wire                CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_counterOnePixelStream_payload;
  reg                 CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_2;
  reg                 CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_counterOnePixelStream_payload_1;
  wire                readStage_counterOnePixelStream_valid;
  wire                readStage_counterOnePixelStream_ready;
  wire       [7:0]    readStage_counterOnePixelStream_payload;
  reg                 CICC1851_readStage_counterOnePixelStream_valid;
  reg        [7:0]    CICC1851_readStage_counterOnePixelStream_payload_2;
  wire                when_Stream_l368_4;
  wire                mainAddrTwoStream_s2mPipe_valid;
  reg                 mainAddrTwoStream_s2mPipe_ready;
  wire       [10:0]   mainAddrTwoStream_s2mPipe_payload;
  reg                 mainAddrTwoStream_rValid;
  reg        [10:0]   mainAddrTwoStream_rData;
  wire                mainAddrTwoStream_s2mPipe_m2sPipe_valid;
  wire                mainAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire       [10:0]   mainAddrTwoStream_s2mPipe_m2sPipe_payload;
  reg                 mainAddrTwoStream_s2mPipe_rValid;
  reg        [10:0]   mainAddrTwoStream_s2mPipe_rData;
  wire                when_Stream_l368_5;
  wire                CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_mainTwoPixelStream_payload;
  reg                 CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_3;
  reg                 CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_mainTwoPixelStream_payload_1;
  wire                readStage_mainTwoPixelStream_valid;
  wire                readStage_mainTwoPixelStream_ready;
  wire       [7:0]    readStage_mainTwoPixelStream_payload;
  reg                 CICC1851_readStage_mainTwoPixelStream_valid;
  reg        [7:0]    CICC1851_readStage_mainTwoPixelStream_payload_2;
  wire                when_Stream_l368_6;
  wire                counterAddrTwoStream_s2mPipe_valid;
  reg                 counterAddrTwoStream_s2mPipe_ready;
  wire       [10:0]   counterAddrTwoStream_s2mPipe_payload;
  reg                 counterAddrTwoStream_rValid;
  reg        [10:0]   counterAddrTwoStream_rData;
  wire                counterAddrTwoStream_s2mPipe_m2sPipe_valid;
  wire                counterAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire       [10:0]   counterAddrTwoStream_s2mPipe_m2sPipe_payload;
  reg                 counterAddrTwoStream_s2mPipe_rValid;
  reg        [10:0]   counterAddrTwoStream_s2mPipe_rData;
  wire                when_Stream_l368_7;
  wire                CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_counterTwoPixelStream_payload;
  reg                 CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_4;
  reg                 CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_counterTwoPixelStream_payload_1;
  wire                readStage_counterTwoPixelStream_valid;
  wire                readStage_counterTwoPixelStream_ready;
  wire       [7:0]    readStage_counterTwoPixelStream_payload;
  reg                 CICC1851_readStage_counterTwoPixelStream_valid;
  reg        [7:0]    CICC1851_readStage_counterTwoPixelStream_payload_2;
  wire                when_Stream_l368_8;
  wire                oddAddrStream_s2mPipe_valid;
  reg                 oddAddrStream_s2mPipe_ready;
  wire       [10:0]   oddAddrStream_s2mPipe_payload;
  reg                 oddAddrStream_rValid;
  reg        [10:0]   oddAddrStream_rData;
  wire                oddAddrStream_s2mPipe_m2sPipe_valid;
  wire                oddAddrStream_s2mPipe_m2sPipe_ready;
  wire       [10:0]   oddAddrStream_s2mPipe_m2sPipe_payload;
  reg                 oddAddrStream_s2mPipe_rValid;
  reg        [10:0]   oddAddrStream_s2mPipe_rData;
  wire                when_Stream_l368_9;
  wire                CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_oddRowPixelStream_payload;
  reg                 CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_5;
  reg                 CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_oddRowPixelStream_payload_1;
  wire                readStage_oddRowPixelStream_valid;
  wire                readStage_oddRowPixelStream_ready;
  wire       [7:0]    readStage_oddRowPixelStream_payload;
  reg                 CICC1851_readStage_oddRowPixelStream_valid;
  reg        [7:0]    CICC1851_readStage_oddRowPixelStream_payload_2;
  wire                when_Stream_l368_10;
  wire                controlStream_s2mPipe_valid;
  reg                 controlStream_s2mPipe_ready;
  wire                controlStream_s2mPipe_payload_frameStart;
  wire                controlStream_s2mPipe_payload_rowEnd;
  wire                controlStream_s2mPipe_payload_passMode;
  wire                controlStream_s2mPipe_payload_passValid;
  wire       [2:0]    controlStream_s2mPipe_payload_onceMode;
  wire                controlStream_s2mPipe_payload_onceValid;
  wire                controlStream_s2mPipe_payload_mainCompare;
  wire                controlStream_s2mPipe_payload_counterCompare;
  wire       [7:0]    controlStream_s2mPipe_payload_mainDiff;
  wire       [7:0]    controlStream_s2mPipe_payload_counterDiff;
  wire                controlStream_s2mPipe_payload_twiceCompValid;
  wire       [2:0]    controlStream_s2mPipe_payload_twiceMode;
  wire                controlStream_s2mPipe_payload_inpValidFlag;
  wire                controlStream_s2mPipe_payload_oddValid;
  reg                 controlStream_rValid;
  reg                 controlStream_rData_frameStart;
  reg                 controlStream_rData_rowEnd;
  reg                 controlStream_rData_passMode;
  reg                 controlStream_rData_passValid;
  reg        [2:0]    controlStream_rData_onceMode;
  reg                 controlStream_rData_onceValid;
  reg                 controlStream_rData_mainCompare;
  reg                 controlStream_rData_counterCompare;
  reg        [7:0]    controlStream_rData_mainDiff;
  reg        [7:0]    controlStream_rData_counterDiff;
  reg                 controlStream_rData_twiceCompValid;
  reg        [2:0]    controlStream_rData_twiceMode;
  reg                 controlStream_rData_inpValidFlag;
  reg                 controlStream_rData_oddValid;
  wire                controlStream_s2mPipe_m2sPipe_valid;
  reg                 controlStream_s2mPipe_m2sPipe_ready;
  wire                controlStream_s2mPipe_m2sPipe_payload_frameStart;
  wire                controlStream_s2mPipe_m2sPipe_payload_rowEnd;
  wire                controlStream_s2mPipe_m2sPipe_payload_passMode;
  wire                controlStream_s2mPipe_m2sPipe_payload_passValid;
  wire       [2:0]    controlStream_s2mPipe_m2sPipe_payload_onceMode;
  wire                controlStream_s2mPipe_m2sPipe_payload_onceValid;
  wire                controlStream_s2mPipe_m2sPipe_payload_mainCompare;
  wire                controlStream_s2mPipe_m2sPipe_payload_counterCompare;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_payload_mainDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_payload_counterDiff;
  wire                controlStream_s2mPipe_m2sPipe_payload_twiceCompValid;
  wire       [2:0]    controlStream_s2mPipe_m2sPipe_payload_twiceMode;
  wire                controlStream_s2mPipe_m2sPipe_payload_inpValidFlag;
  wire                controlStream_s2mPipe_m2sPipe_payload_oddValid;
  reg                 controlStream_s2mPipe_rValid;
  reg                 controlStream_s2mPipe_rData_frameStart;
  reg                 controlStream_s2mPipe_rData_rowEnd;
  reg                 controlStream_s2mPipe_rData_passMode;
  reg                 controlStream_s2mPipe_rData_passValid;
  reg        [2:0]    controlStream_s2mPipe_rData_onceMode;
  reg                 controlStream_s2mPipe_rData_onceValid;
  reg                 controlStream_s2mPipe_rData_mainCompare;
  reg                 controlStream_s2mPipe_rData_counterCompare;
  reg        [7:0]    controlStream_s2mPipe_rData_mainDiff;
  reg        [7:0]    controlStream_s2mPipe_rData_counterDiff;
  reg                 controlStream_s2mPipe_rData_twiceCompValid;
  reg        [2:0]    controlStream_s2mPipe_rData_twiceMode;
  reg                 controlStream_s2mPipe_rData_inpValidFlag;
  reg                 controlStream_s2mPipe_rData_oddValid;
  wire                when_Stream_l368_11;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_valid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_ready;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_frameStart;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_rowEnd;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passMode;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passValid;
  wire       [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceMode;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceValid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainCompare;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterCompare;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDiff;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceCompValid;
  wire       [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceMode;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_inpValidFlag;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_oddValid;
  reg                 controlStream_s2mPipe_m2sPipe_rValid;
  reg                 controlStream_s2mPipe_m2sPipe_rData_frameStart;
  reg                 controlStream_s2mPipe_m2sPipe_rData_rowEnd;
  reg                 controlStream_s2mPipe_m2sPipe_rData_passMode;
  reg                 controlStream_s2mPipe_m2sPipe_rData_passValid;
  reg        [2:0]    controlStream_s2mPipe_m2sPipe_rData_onceMode;
  reg                 controlStream_s2mPipe_m2sPipe_rData_onceValid;
  reg                 controlStream_s2mPipe_m2sPipe_rData_mainCompare;
  reg                 controlStream_s2mPipe_m2sPipe_rData_counterCompare;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_rData_mainDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_rData_counterDiff;
  reg                 controlStream_s2mPipe_m2sPipe_rData_twiceCompValid;
  reg        [2:0]    controlStream_s2mPipe_m2sPipe_rData_twiceMode;
  reg                 controlStream_s2mPipe_m2sPipe_rData_inpValidFlag;
  reg                 controlStream_s2mPipe_m2sPipe_rData_oddValid;
  wire                when_Stream_l368_12;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_valid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_frameStart;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_rowEnd;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_passMode;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_passValid;
  wire       [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_onceMode;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_onceValid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainCompare;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterCompare;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterDiff;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_twiceCompValid;
  wire       [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_twiceMode;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_inpValidFlag;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_oddValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_frameStart;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_rowEnd;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_passMode;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_passValid;
  reg        [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_onceMode;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_onceValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainCompare;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterCompare;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterDiff;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_twiceCompValid;
  reg        [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_twiceMode;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_inpValidFlag;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_oddValid;
  wire                readStage_controlPipe_valid;
  wire                readStage_controlPipe_ready;
  wire                readStage_controlPipe_payload_frameStart;
  wire                readStage_controlPipe_payload_rowEnd;
  wire                readStage_controlPipe_payload_passMode;
  wire                readStage_controlPipe_payload_passValid;
  wire       [2:0]    readStage_controlPipe_payload_onceMode;
  wire                readStage_controlPipe_payload_onceValid;
  wire                readStage_controlPipe_payload_mainCompare;
  wire                readStage_controlPipe_payload_counterCompare;
  wire       [7:0]    readStage_controlPipe_payload_mainDiff;
  wire       [7:0]    readStage_controlPipe_payload_counterDiff;
  wire                readStage_controlPipe_payload_twiceCompValid;
  wire       [2:0]    readStage_controlPipe_payload_twiceMode;
  wire                readStage_controlPipe_payload_inpValidFlag;
  wire                readStage_controlPipe_payload_oddValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_frameStart;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_rowEnd;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_passMode;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_passValid;
  reg        [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_onceMode;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_onceValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainCompare;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterCompare;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterDiff;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_twiceCompValid;
  reg        [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_twiceMode;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_inpValidFlag;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_oddValid;
  wire                when_Stream_l368_13;
  wire                readStage_mainOnePixelStream_s2mPipe_valid;
  reg                 readStage_mainOnePixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_mainOnePixelStream_s2mPipe_payload;
  reg                 readStage_mainOnePixelStream_rValid;
  reg        [7:0]    readStage_mainOnePixelStream_rData;
  wire                compareStage_mainOnePixelStream_valid;
  wire                compareStage_mainOnePixelStream_ready;
  wire       [7:0]    compareStage_mainOnePixelStream_payload;
  reg                 readStage_mainOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_mainOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_14;
  wire                readStage_counterOnePixelStream_s2mPipe_valid;
  reg                 readStage_counterOnePixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_counterOnePixelStream_s2mPipe_payload;
  reg                 readStage_counterOnePixelStream_rValid;
  reg        [7:0]    readStage_counterOnePixelStream_rData;
  wire                compareStage_counterOnePixelStream_valid;
  wire                compareStage_counterOnePixelStream_ready;
  wire       [7:0]    compareStage_counterOnePixelStream_payload;
  reg                 readStage_counterOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_counterOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_15;
  wire                readStage_mainTwoPixelStream_s2mPipe_valid;
  reg                 readStage_mainTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_mainTwoPixelStream_s2mPipe_payload;
  reg                 readStage_mainTwoPixelStream_rValid;
  reg        [7:0]    readStage_mainTwoPixelStream_rData;
  wire                compareStage_mainTwoPixelStream_valid;
  wire                compareStage_mainTwoPixelStream_ready;
  wire       [7:0]    compareStage_mainTwoPixelStream_payload;
  reg                 readStage_mainTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_mainTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_16;
  wire                readStage_counterTwoPixelStream_s2mPipe_valid;
  reg                 readStage_counterTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_counterTwoPixelStream_s2mPipe_payload;
  reg                 readStage_counterTwoPixelStream_rValid;
  reg        [7:0]    readStage_counterTwoPixelStream_rData;
  wire                compareStage_counterTwoPixelStream_valid;
  wire                compareStage_counterTwoPixelStream_ready;
  wire       [7:0]    compareStage_counterTwoPixelStream_payload;
  reg                 readStage_counterTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_counterTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_17;
  wire                readStage_oddRowPixelStream_s2mPipe_valid;
  reg                 readStage_oddRowPixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_oddRowPixelStream_s2mPipe_payload;
  reg                 readStage_oddRowPixelStream_rValid;
  reg        [7:0]    readStage_oddRowPixelStream_rData;
  wire                compareStage_oddRowPixelStream_valid;
  wire                compareStage_oddRowPixelStream_ready;
  wire       [7:0]    compareStage_oddRowPixelStream_payload;
  reg                 readStage_oddRowPixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_oddRowPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_18;
  reg                 CICC1851_readStage_controlPipe_translated_payload_mainCompare;
  reg                 CICC1851_readStage_controlPipe_translated_payload_counterCompare;
  wire                when_SuperResolutionPart2_l290;
  wire                when_SuperResolutionPart2_l294;
  wire                when_SuperResolutionPart2_l298;
  wire                when_SuperResolutionPart2_l302;
  wire                when_SuperResolutionPart2_l313;
  wire                when_SuperResolutionPart2_l315;
  wire                when_SuperResolutionPart2_l319;
  wire                when_SuperResolutionPart2_l321;
  wire                when_SuperResolutionPart2_l326;
  wire                when_SuperResolutionPart2_l331;
  wire                readStage_controlPipe_translated_valid;
  wire                readStage_controlPipe_translated_ready;
  wire                readStage_controlPipe_translated_payload_frameStart;
  wire                readStage_controlPipe_translated_payload_rowEnd;
  wire                readStage_controlPipe_translated_payload_passMode;
  wire                readStage_controlPipe_translated_payload_passValid;
  wire       [2:0]    readStage_controlPipe_translated_payload_onceMode;
  wire                readStage_controlPipe_translated_payload_onceValid;
  wire                readStage_controlPipe_translated_payload_mainCompare;
  wire                readStage_controlPipe_translated_payload_counterCompare;
  wire       [7:0]    readStage_controlPipe_translated_payload_mainDiff;
  wire       [7:0]    readStage_controlPipe_translated_payload_counterDiff;
  wire                readStage_controlPipe_translated_payload_twiceCompValid;
  wire       [2:0]    readStage_controlPipe_translated_payload_twiceMode;
  wire                readStage_controlPipe_translated_payload_inpValidFlag;
  wire                readStage_controlPipe_translated_payload_oddValid;
  wire                readStage_controlPipe_translated_s2mPipe_valid;
  reg                 readStage_controlPipe_translated_s2mPipe_ready;
  wire                readStage_controlPipe_translated_s2mPipe_payload_frameStart;
  wire                readStage_controlPipe_translated_s2mPipe_payload_rowEnd;
  wire                readStage_controlPipe_translated_s2mPipe_payload_passMode;
  wire                readStage_controlPipe_translated_s2mPipe_payload_passValid;
  wire       [2:0]    readStage_controlPipe_translated_s2mPipe_payload_onceMode;
  wire                readStage_controlPipe_translated_s2mPipe_payload_onceValid;
  wire                readStage_controlPipe_translated_s2mPipe_payload_mainCompare;
  wire                readStage_controlPipe_translated_s2mPipe_payload_counterCompare;
  wire       [7:0]    readStage_controlPipe_translated_s2mPipe_payload_mainDiff;
  wire       [7:0]    readStage_controlPipe_translated_s2mPipe_payload_counterDiff;
  wire                readStage_controlPipe_translated_s2mPipe_payload_twiceCompValid;
  wire       [2:0]    readStage_controlPipe_translated_s2mPipe_payload_twiceMode;
  wire                readStage_controlPipe_translated_s2mPipe_payload_inpValidFlag;
  wire                readStage_controlPipe_translated_s2mPipe_payload_oddValid;
  reg                 readStage_controlPipe_translated_rValid;
  reg                 readStage_controlPipe_translated_rData_frameStart;
  reg                 readStage_controlPipe_translated_rData_rowEnd;
  reg                 readStage_controlPipe_translated_rData_passMode;
  reg                 readStage_controlPipe_translated_rData_passValid;
  reg        [2:0]    readStage_controlPipe_translated_rData_onceMode;
  reg                 readStage_controlPipe_translated_rData_onceValid;
  reg                 readStage_controlPipe_translated_rData_mainCompare;
  reg                 readStage_controlPipe_translated_rData_counterCompare;
  reg        [7:0]    readStage_controlPipe_translated_rData_mainDiff;
  reg        [7:0]    readStage_controlPipe_translated_rData_counterDiff;
  reg                 readStage_controlPipe_translated_rData_twiceCompValid;
  reg        [2:0]    readStage_controlPipe_translated_rData_twiceMode;
  reg                 readStage_controlPipe_translated_rData_inpValidFlag;
  reg                 readStage_controlPipe_translated_rData_oddValid;
  wire                compareStage_controlPipe_valid;
  wire                compareStage_controlPipe_ready;
  wire                compareStage_controlPipe_payload_frameStart;
  wire                compareStage_controlPipe_payload_rowEnd;
  wire                compareStage_controlPipe_payload_passMode;
  wire                compareStage_controlPipe_payload_passValid;
  wire       [2:0]    compareStage_controlPipe_payload_onceMode;
  wire                compareStage_controlPipe_payload_onceValid;
  wire                compareStage_controlPipe_payload_mainCompare;
  wire                compareStage_controlPipe_payload_counterCompare;
  wire       [7:0]    compareStage_controlPipe_payload_mainDiff;
  wire       [7:0]    compareStage_controlPipe_payload_counterDiff;
  wire                compareStage_controlPipe_payload_twiceCompValid;
  wire       [2:0]    compareStage_controlPipe_payload_twiceMode;
  wire                compareStage_controlPipe_payload_inpValidFlag;
  wire                compareStage_controlPipe_payload_oddValid;
  reg                 readStage_controlPipe_translated_s2mPipe_rValid;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_frameStart;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_rowEnd;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_passMode;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_passValid;
  reg        [2:0]    readStage_controlPipe_translated_s2mPipe_rData_onceMode;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_onceValid;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_mainCompare;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_counterCompare;
  reg        [7:0]    readStage_controlPipe_translated_s2mPipe_rData_mainDiff;
  reg        [7:0]    readStage_controlPipe_translated_s2mPipe_rData_counterDiff;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_twiceCompValid;
  reg        [2:0]    readStage_controlPipe_translated_s2mPipe_rData_twiceMode;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_inpValidFlag;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_oddValid;
  wire                when_Stream_l368_19;
  wire                compareStage_mainOnePixelStream_s2mPipe_valid;
  reg                 compareStage_mainOnePixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_mainOnePixelStream_s2mPipe_payload;
  reg                 compareStage_mainOnePixelStream_rValid;
  reg        [7:0]    compareStage_mainOnePixelStream_rData;
  wire                diffStage_mainOnePixelStream_valid;
  wire                diffStage_mainOnePixelStream_ready;
  wire       [7:0]    diffStage_mainOnePixelStream_payload;
  reg                 compareStage_mainOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_mainOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_20;
  wire                compareStage_counterOnePixelStream_s2mPipe_valid;
  reg                 compareStage_counterOnePixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_counterOnePixelStream_s2mPipe_payload;
  reg                 compareStage_counterOnePixelStream_rValid;
  reg        [7:0]    compareStage_counterOnePixelStream_rData;
  wire                diffStage_counterOnePixelStream_valid;
  wire                diffStage_counterOnePixelStream_ready;
  wire       [7:0]    diffStage_counterOnePixelStream_payload;
  reg                 compareStage_counterOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_counterOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_21;
  wire                compareStage_mainTwoPixelStream_s2mPipe_valid;
  reg                 compareStage_mainTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_mainTwoPixelStream_s2mPipe_payload;
  reg                 compareStage_mainTwoPixelStream_rValid;
  reg        [7:0]    compareStage_mainTwoPixelStream_rData;
  wire                diffStage_mainTwoPixelStream_valid;
  wire                diffStage_mainTwoPixelStream_ready;
  wire       [7:0]    diffStage_mainTwoPixelStream_payload;
  reg                 compareStage_mainTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_mainTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_22;
  wire                compareStage_counterTwoPixelStream_s2mPipe_valid;
  reg                 compareStage_counterTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_counterTwoPixelStream_s2mPipe_payload;
  reg                 compareStage_counterTwoPixelStream_rValid;
  reg        [7:0]    compareStage_counterTwoPixelStream_rData;
  wire                diffStage_counterTwoPixelStream_valid;
  wire                diffStage_counterTwoPixelStream_ready;
  wire       [7:0]    diffStage_counterTwoPixelStream_payload;
  reg                 compareStage_counterTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_counterTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_23;
  wire                compareStage_oddRowPixelStream_s2mPipe_valid;
  reg                 compareStage_oddRowPixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_oddRowPixelStream_s2mPipe_payload;
  reg                 compareStage_oddRowPixelStream_rValid;
  reg        [7:0]    compareStage_oddRowPixelStream_rData;
  wire                diffStage_oddRowPixelStream_valid;
  wire                diffStage_oddRowPixelStream_ready;
  wire       [7:0]    diffStage_oddRowPixelStream_payload;
  reg                 compareStage_oddRowPixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_oddRowPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_24;
  reg        [7:0]    CICC1851_compareStage_controlPipe_translated_payload_mainDiff;
  reg        [7:0]    CICC1851_compareStage_controlPipe_translated_payload_counterDiff;
  wire                compareStage_controlPipe_translated_valid;
  wire                compareStage_controlPipe_translated_ready;
  wire                compareStage_controlPipe_translated_payload_frameStart;
  wire                compareStage_controlPipe_translated_payload_rowEnd;
  wire                compareStage_controlPipe_translated_payload_passMode;
  wire                compareStage_controlPipe_translated_payload_passValid;
  wire       [2:0]    compareStage_controlPipe_translated_payload_onceMode;
  wire                compareStage_controlPipe_translated_payload_onceValid;
  wire                compareStage_controlPipe_translated_payload_mainCompare;
  wire                compareStage_controlPipe_translated_payload_counterCompare;
  wire       [7:0]    compareStage_controlPipe_translated_payload_mainDiff;
  wire       [7:0]    compareStage_controlPipe_translated_payload_counterDiff;
  wire                compareStage_controlPipe_translated_payload_twiceCompValid;
  wire       [2:0]    compareStage_controlPipe_translated_payload_twiceMode;
  wire                compareStage_controlPipe_translated_payload_inpValidFlag;
  wire                compareStage_controlPipe_translated_payload_oddValid;
  wire                compareStage_controlPipe_translated_s2mPipe_valid;
  reg                 compareStage_controlPipe_translated_s2mPipe_ready;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_frameStart;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_rowEnd;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_passMode;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_passValid;
  wire       [2:0]    compareStage_controlPipe_translated_s2mPipe_payload_onceMode;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_onceValid;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_mainCompare;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_counterCompare;
  wire       [7:0]    compareStage_controlPipe_translated_s2mPipe_payload_mainDiff;
  wire       [7:0]    compareStage_controlPipe_translated_s2mPipe_payload_counterDiff;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_twiceCompValid;
  wire       [2:0]    compareStage_controlPipe_translated_s2mPipe_payload_twiceMode;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_inpValidFlag;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_oddValid;
  reg                 compareStage_controlPipe_translated_rValid;
  reg                 compareStage_controlPipe_translated_rData_frameStart;
  reg                 compareStage_controlPipe_translated_rData_rowEnd;
  reg                 compareStage_controlPipe_translated_rData_passMode;
  reg                 compareStage_controlPipe_translated_rData_passValid;
  reg        [2:0]    compareStage_controlPipe_translated_rData_onceMode;
  reg                 compareStage_controlPipe_translated_rData_onceValid;
  reg                 compareStage_controlPipe_translated_rData_mainCompare;
  reg                 compareStage_controlPipe_translated_rData_counterCompare;
  reg        [7:0]    compareStage_controlPipe_translated_rData_mainDiff;
  reg        [7:0]    compareStage_controlPipe_translated_rData_counterDiff;
  reg                 compareStage_controlPipe_translated_rData_twiceCompValid;
  reg        [2:0]    compareStage_controlPipe_translated_rData_twiceMode;
  reg                 compareStage_controlPipe_translated_rData_inpValidFlag;
  reg                 compareStage_controlPipe_translated_rData_oddValid;
  wire                diffStage_controlPipe_valid;
  wire                diffStage_controlPipe_ready;
  wire                diffStage_controlPipe_payload_frameStart;
  wire                diffStage_controlPipe_payload_rowEnd;
  wire                diffStage_controlPipe_payload_passMode;
  wire                diffStage_controlPipe_payload_passValid;
  wire       [2:0]    diffStage_controlPipe_payload_onceMode;
  wire                diffStage_controlPipe_payload_onceValid;
  wire                diffStage_controlPipe_payload_mainCompare;
  wire                diffStage_controlPipe_payload_counterCompare;
  wire       [7:0]    diffStage_controlPipe_payload_mainDiff;
  wire       [7:0]    diffStage_controlPipe_payload_counterDiff;
  wire                diffStage_controlPipe_payload_twiceCompValid;
  wire       [2:0]    diffStage_controlPipe_payload_twiceMode;
  wire                diffStage_controlPipe_payload_inpValidFlag;
  wire                diffStage_controlPipe_payload_oddValid;
  reg                 compareStage_controlPipe_translated_s2mPipe_rValid;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_frameStart;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_rowEnd;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_passMode;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_passValid;
  reg        [2:0]    compareStage_controlPipe_translated_s2mPipe_rData_onceMode;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_onceValid;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_mainCompare;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_counterCompare;
  reg        [7:0]    compareStage_controlPipe_translated_s2mPipe_rData_mainDiff;
  reg        [7:0]    compareStage_controlPipe_translated_s2mPipe_rData_counterDiff;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_twiceCompValid;
  reg        [2:0]    compareStage_controlPipe_translated_s2mPipe_rData_twiceMode;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_inpValidFlag;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_oddValid;
  wire                when_Stream_l368_25;
  wire                diffStage_mainOnePixelStream_s2mPipe_valid;
  reg                 diffStage_mainOnePixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_mainOnePixelStream_s2mPipe_payload;
  reg                 diffStage_mainOnePixelStream_rValid;
  reg        [7:0]    diffStage_mainOnePixelStream_rData;
  wire                resultStage_mainOnePixelStream_valid;
  wire                resultStage_mainOnePixelStream_ready;
  wire       [7:0]    resultStage_mainOnePixelStream_payload;
  reg                 diffStage_mainOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_mainOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_26;
  wire                diffStage_counterOnePixelStream_s2mPipe_valid;
  reg                 diffStage_counterOnePixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_counterOnePixelStream_s2mPipe_payload;
  reg                 diffStage_counterOnePixelStream_rValid;
  reg        [7:0]    diffStage_counterOnePixelStream_rData;
  wire                resultStage_counterOnePixelStream_valid;
  wire                resultStage_counterOnePixelStream_ready;
  wire       [7:0]    resultStage_counterOnePixelStream_payload;
  reg                 diffStage_counterOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_counterOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_27;
  wire                diffStage_mainTwoPixelStream_s2mPipe_valid;
  reg                 diffStage_mainTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_mainTwoPixelStream_s2mPipe_payload;
  reg                 diffStage_mainTwoPixelStream_rValid;
  reg        [7:0]    diffStage_mainTwoPixelStream_rData;
  wire                resultStage_mainTwoPixelStream_valid;
  wire                resultStage_mainTwoPixelStream_ready;
  wire       [7:0]    resultStage_mainTwoPixelStream_payload;
  reg                 diffStage_mainTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_mainTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_28;
  wire                diffStage_counterTwoPixelStream_s2mPipe_valid;
  reg                 diffStage_counterTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_counterTwoPixelStream_s2mPipe_payload;
  reg                 diffStage_counterTwoPixelStream_rValid;
  reg        [7:0]    diffStage_counterTwoPixelStream_rData;
  wire                resultStage_counterTwoPixelStream_valid;
  wire                resultStage_counterTwoPixelStream_ready;
  wire       [7:0]    resultStage_counterTwoPixelStream_payload;
  reg                 diffStage_counterTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_counterTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_29;
  wire                diffStage_oddRowPixelStream_s2mPipe_valid;
  reg                 diffStage_oddRowPixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_oddRowPixelStream_s2mPipe_payload;
  reg                 diffStage_oddRowPixelStream_rValid;
  reg        [7:0]    diffStage_oddRowPixelStream_rData;
  wire                resultStage_oddRowPixelStream_valid;
  wire                resultStage_oddRowPixelStream_ready;
  wire       [7:0]    resultStage_oddRowPixelStream_payload;
  reg                 diffStage_oddRowPixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_oddRowPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_30;
  wire       [2:0]    CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceMode;
  wire                CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceValid;
  wire       [7:0]    CICC1851_when_SuperResolutionPart2_l419;
  wire       [7:0]    CICC1851_when_SuperResolutionPart2_l428;
  wire                CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceCompValid;
  wire       [2:0]    CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceMode;
  reg                 CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag;
  wire                when_SuperResolutionPart2_l419;
  wire                when_SuperResolutionPart2_l420;
  wire                when_SuperResolutionPart2_l421;
  wire                when_SuperResolutionPart2_l422;
  wire                when_SuperResolutionPart2_l428;
  wire                when_SuperResolutionPart2_l429;
  wire                when_SuperResolutionPart2_l430;
  wire                when_SuperResolutionPart2_l431;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_valid;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_ready;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_payload_frameStart;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_payload_rowEnd;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_payload_passMode;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_payload_passValid;
  wire       [2:0]    diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceMode;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceValid;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_payload_mainCompare;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_payload_counterCompare;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_translated_payload_mainDiff;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_translated_payload_counterDiff;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceCompValid;
  wire       [2:0]    diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceMode;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_payload_oddValid;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_valid;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_ready;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_frameStart;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_rowEnd;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_passMode;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_passValid;
  wire       [2:0]    diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_onceMode;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_onceValid;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_mainCompare;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_counterCompare;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_mainDiff;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_counterDiff;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_twiceCompValid;
  wire       [2:0]    diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_twiceMode;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_inpValidFlag;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_oddValid;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_rValid;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_rData_frameStart;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_rData_rowEnd;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_rData_passMode;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_rData_passValid;
  reg        [2:0]    diffStage_controlPipe_fork_io_outputs_0_translated_rData_onceMode;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_rData_onceValid;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_rData_mainCompare;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_rData_counterCompare;
  reg        [7:0]    diffStage_controlPipe_fork_io_outputs_0_translated_rData_mainDiff;
  reg        [7:0]    diffStage_controlPipe_fork_io_outputs_0_translated_rData_counterDiff;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_rData_twiceCompValid;
  reg        [2:0]    diffStage_controlPipe_fork_io_outputs_0_translated_rData_twiceMode;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_rData_inpValidFlag;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_rData_oddValid;
  wire                resultStage_controlPipe_valid;
  wire                resultStage_controlPipe_ready;
  wire                resultStage_controlPipe_payload_frameStart;
  wire                resultStage_controlPipe_payload_rowEnd;
  wire                resultStage_controlPipe_payload_passMode;
  wire                resultStage_controlPipe_payload_passValid;
  wire       [2:0]    resultStage_controlPipe_payload_onceMode;
  wire                resultStage_controlPipe_payload_onceValid;
  wire                resultStage_controlPipe_payload_mainCompare;
  wire                resultStage_controlPipe_payload_counterCompare;
  wire       [7:0]    resultStage_controlPipe_payload_mainDiff;
  wire       [7:0]    resultStage_controlPipe_payload_counterDiff;
  wire                resultStage_controlPipe_payload_twiceCompValid;
  wire       [2:0]    resultStage_controlPipe_payload_twiceMode;
  wire                resultStage_controlPipe_payload_inpValidFlag;
  wire                resultStage_controlPipe_payload_oddValid;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rValid;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_frameStart;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_rowEnd;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_passMode;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_passValid;
  reg        [2:0]    diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_onceMode;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_onceValid;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_mainCompare;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_counterCompare;
  reg        [7:0]    diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_mainDiff;
  reg        [7:0]    diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_counterDiff;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_twiceCompValid;
  reg        [2:0]    diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_twiceMode;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_inpValidFlag;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_oddValid;
  wire                when_Stream_l368_31;
  wire                resultStage_pixelStream_valid;
  wire                resultStage_pixelStream_ready;
  reg        [7:0]    resultStage_pixelStream_payload;
  wire                when_SuperResolutionPart2_l451;
  wire                when_SuperResolutionPart2_l455;
  wire                when_SuperResolutionPart2_l459;
  wire                when_SuperResolutionPart2_l463;
  wire                when_SuperResolutionPart2_l474;
  wire                when_SuperResolutionPart2_l477;
  wire                when_SuperResolutionPart2_l482;
  wire                when_SuperResolutionPart2_l485;
  wire                when_SuperResolutionPart2_l491;
  wire                when_SuperResolutionPart2_l496;
  wire                resultStage_pixelStream_s2mPipe_valid;
  reg                 resultStage_pixelStream_s2mPipe_ready;
  wire       [7:0]    resultStage_pixelStream_s2mPipe_payload;
  reg                 resultStage_pixelStream_rValid;
  reg        [7:0]    resultStage_pixelStream_rData;
  wire                resultStage_resultStream_valid;
  wire                resultStage_resultStream_ready;
  wire       [7:0]    resultStage_resultStream_payload;
  reg                 resultStage_pixelStream_s2mPipe_rValid;
  reg        [7:0]    resultStage_pixelStream_s2mPipe_rData;
  wire                when_Stream_l368_32;
  wire                CICC1851_resultStage_mainOnePixelStream_ready;
  reg                 CICC1851_resultStage_mainOnePixelStream_ready_1;
  wire                CICC1851_resultStage_mainOnePixelStream_ready_2;
  wire                when_Stream_l438;
  reg                 resultsJoin_valid;
  wire                resultsJoin_ready;
  wire                pixelsStream_valid;
  wire                pixelsStream_ready;
  wire       [7:0]    pixelsStream_payload_pixel;
  wire                pixelsStream_payload_frameStart;
  wire                pixelsStream_payload_rowEnd;
  wire                pixelsStream_payload_inpValid;
  wire                pixelsStream_s2mPipe_valid;
  reg                 pixelsStream_s2mPipe_ready;
  wire       [7:0]    pixelsStream_s2mPipe_payload_pixel;
  wire                pixelsStream_s2mPipe_payload_frameStart;
  wire                pixelsStream_s2mPipe_payload_rowEnd;
  wire                pixelsStream_s2mPipe_payload_inpValid;
  reg                 pixelsStream_rValid;
  reg        [7:0]    pixelsStream_rData_pixel;
  reg                 pixelsStream_rData_frameStart;
  reg                 pixelsStream_rData_rowEnd;
  reg                 pixelsStream_rData_inpValid;
  wire                pixelsStream_s2mPipe_m2sPipe_valid;
  wire                pixelsStream_s2mPipe_m2sPipe_ready;
  wire       [7:0]    pixelsStream_s2mPipe_m2sPipe_payload_pixel;
  wire                pixelsStream_s2mPipe_m2sPipe_payload_frameStart;
  wire                pixelsStream_s2mPipe_m2sPipe_payload_rowEnd;
  wire                pixelsStream_s2mPipe_m2sPipe_payload_inpValid;
  reg                 pixelsStream_s2mPipe_rValid;
  reg        [7:0]    pixelsStream_s2mPipe_rData_pixel;
  reg                 pixelsStream_s2mPipe_rData_frameStart;
  reg                 pixelsStream_s2mPipe_rData_rowEnd;
  reg                 pixelsStream_s2mPipe_rData_inpValid;
  wire                when_Stream_l368_33;
  wire                controlStateMachine_wantExit;
  reg                 controlStateMachine_wantStart;
  wire                controlStateMachine_wantKill;
  wire                when_SuperResolutionPart2_l761;
  wire                controlStream_fire_4;
  wire                when_SuperResolutionPart2_l763;
  wire                controlStream_fire_5;
  wire                when_SuperResolutionPart2_l764;
  wire                controlStream_fire_6;
  wire                when_SuperResolutionPart2_l766;
  wire                controlStream_fire_7;
  wire                when_SuperResolutionPart2_l783;
  wire                when_SuperResolutionPart2_l785;
  wire                when_SuperResolutionPart2_l787;
  wire                when_SuperResolutionPart2_l789;
  wire                when_SuperResolutionPart2_l793;
  wire                when_SuperResolutionPart2_l796;
  wire                when_SuperResolutionPart2_l799;
  wire                when_SuperResolutionPart2_l802;
  reg        [2:0]    controlStateMachine_stateReg;
  reg        [2:0]    controlStateMachine_stateNext;
  wire                passPixels_fire_13;
  wire                passPixels_fire_14;
  wire                passPixels_fire_15;
  wire                passPixels_fire_16;
  wire                when_SuperResolutionPart2_l560;
  wire                controlStream_fire_8;
  wire                passPixels_fire_17;
  wire                when_SuperResolutionPart2_l573;
  wire                passPixels_fire_18;
  wire                when_SuperResolutionPart2_l578;
  wire                when_SuperResolutionPart2_l585;
  wire                when_SuperResolutionPart2_l588;
  wire                passPixels_fire_19;
  wire                when_SuperResolutionPart2_l590;
  wire                when_SuperResolutionPart2_l602;
  wire                when_SuperResolutionPart2_l603;
  wire                when_SuperResolutionPart2_l605;
  wire                when_SuperResolutionPart2_l606;
  wire                when_SuperResolutionPart2_l609;
  wire                controlStream_fire_9;
  wire                when_SuperResolutionPart2_l630;
  wire                controlStream_fire_10;
  wire                passPixels_fire_20;
  wire                when_SuperResolutionPart2_l642;
  wire                passPixels_fire_21;
  wire                when_SuperResolutionPart2_l647;
  wire                passPixels_fire_22;
  wire                when_SuperResolutionPart2_l653;
  wire                passPixels_fire_23;
  wire                when_SuperResolutionPart2_l662;
  wire                when_SuperResolutionPart2_l667;
  wire                when_SuperResolutionPart2_l668;
  wire                controlStream_fire_11;
  `ifndef SYNTHESIS
  reg [39:0] controlStateMachine_stateReg_string;
  reg [39:0] controlStateMachine_stateNext_string;
  `endif

  reg [7:0] lineBufferOne [0:1919];
  reg [7:0] lineBufferTwo [0:1919];
  reg [7:0] lineBufferOdd [0:1919];

  assign CICC1851_bufferRowCount_valueNext_1 = bufferRowCount_willIncrement;
  assign CICC1851_bufferRowCount_valueNext = {10'd0, CICC1851_bufferRowCount_valueNext_1};
  assign CICC1851_bufferWAddr_valueNext_1 = bufferWAddr_willIncrement;
  assign CICC1851_bufferWAddr_valueNext = {10'd0, CICC1851_bufferWAddr_valueNext_1};
  assign CICC1851_outPixelAddr_valueNext_1 = outPixelAddr_willIncrement;
  assign CICC1851_outPixelAddr_valueNext = {11'd0, CICC1851_outPixelAddr_valueNext_1};
  assign CICC1851_outRowCount_valueNext_1 = outRowCount_willIncrement;
  assign CICC1851_outRowCount_valueNext = {11'd0, CICC1851_outRowCount_valueNext_1};
  assign CICC1851_alreadySendRow_valueNext_1 = alreadySendRow_willIncrement;
  assign CICC1851_alreadySendRow_valueNext = {11'd0, CICC1851_alreadySendRow_valueNext_1};
  assign CICC1851_alreadySendCountInRow_valueNext_1 = alreadySendCountInRow_willIncrement;
  assign CICC1851_alreadySendCountInRow_valueNext = {11'd0, CICC1851_alreadySendCountInRow_valueNext_1};
  assign CICC1851_mainAddrOne = (outPixelAddr_value / 2'b10);
  assign CICC1851_counterAddrOne = (outPixelAddr_value / 2'b10);
  assign CICC1851_mainAddrTwo = (outPixelAddr_value / 2'b10);
  assign CICC1851_counterAddrTwo = (outPixelAddr_value / 2'b10);
  assign CICC1851_oddAddr = (outPixelAddr_value / 2'b10);
  assign CICC1851_when_SuperResolutionPart2_l181 = {1'd0, bufferWAddr_value};
  assign CICC1851_when_SuperResolutionPart2_l181_1 = (CICC1851_when_SuperResolutionPart2_l181_2 - 12'h002);
  assign CICC1851_when_SuperResolutionPart2_l181_2 = (2'b10 * bmpWidth);
  assign CICC1851_when_SuperResolutionPart2_l182 = {1'd0, bufferRowCount_value};
  assign CICC1851_when_SuperResolutionPart2_l182_1 = (CICC1851_when_SuperResolutionPart2_l182_2 - 12'h002);
  assign CICC1851_when_SuperResolutionPart2_l182_2 = (2'b10 * bmpHeight);
  assign CICC1851_when_SuperResolutionPart2_l195 = (bufferRowCount_value % 2'b10);
  assign CICC1851_when_SuperResolutionPart2_l218 = (outRowCount_value % 3'b100);
  assign CICC1851_when_SuperResolutionPart2_l234 = {1'd0, alreadySendCountInRow_value};
  assign CICC1851_when_SuperResolutionPart2_l234_1 = (CICC1851_when_SuperResolutionPart2_l234_2 - 13'h0002);
  assign CICC1851_when_SuperResolutionPart2_l234_2 = (3'b100 * bmpWidth);
  assign CICC1851_when_SuperResolutionPart2_l235 = {1'd0, alreadySendRow_value};
  assign CICC1851_when_SuperResolutionPart2_l235_1 = (CICC1851_when_SuperResolutionPart2_l235_2 - 13'h0002);
  assign CICC1851_when_SuperResolutionPart2_l235_2 = (3'b100 * bmpHeight);
  assign CICC1851_resultStage_pixelStream_payload = (CICC1851_resultStage_pixelStream_payload_1 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_1 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_2 = (CICC1851_resultStage_pixelStream_payload_3 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_3 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_4 = (CICC1851_resultStage_pixelStream_payload_5 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_5 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_mainTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_6 = (CICC1851_resultStage_pixelStream_payload_7 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_7 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_mainOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_8 = (CICC1851_resultStage_pixelStream_payload_9 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_9 = ({1'b0,diffStage_counterOnePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_10 = (CICC1851_resultStage_pixelStream_payload_11 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_11 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_mainTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_12 = (CICC1851_resultStage_pixelStream_payload_13 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_13 = ({1'b0,diffStage_counterOnePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_14 = (CICC1851_resultStage_pixelStream_payload_15 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_15 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_mainTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_16 = (CICC1851_resultStage_pixelStream_payload_17 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_17 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_18 = (CICC1851_resultStage_pixelStream_payload_19 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_19 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_when_SuperResolutionPart2_l763 = {1'd0, outPixelAddr_value};
  assign CICC1851_when_SuperResolutionPart2_l763_1 = (CICC1851_when_SuperResolutionPart2_l763_2 - 13'h0002);
  assign CICC1851_when_SuperResolutionPart2_l763_2 = (3'b100 * bmpWidth);
  assign CICC1851_when_SuperResolutionPart2_l764 = {1'd0, outRowCount_value};
  assign CICC1851_when_SuperResolutionPart2_l764_1 = (CICC1851_when_SuperResolutionPart2_l764_2 - 13'h0002);
  assign CICC1851_when_SuperResolutionPart2_l764_2 = (3'b100 * bmpHeight);
  assign CICC1851_when_SuperResolutionPart2_l783 = (outRowCount_value % 3'b100);
  assign CICC1851_when_SuperResolutionPart2_l785 = (outRowCount_value % 3'b100);
  assign CICC1851_when_SuperResolutionPart2_l787 = (outRowCount_value % 3'b100);
  assign CICC1851_when_SuperResolutionPart2_l789 = (outRowCount_value % 3'b100);
  assign CICC1851_when_SuperResolutionPart2_l793 = (outPixelAddr_value % 3'b100);
  assign CICC1851_when_SuperResolutionPart2_l796 = (outPixelAddr_value % 3'b100);
  assign CICC1851_when_SuperResolutionPart2_l799 = (outPixelAddr_value % 3'b100);
  assign CICC1851_when_SuperResolutionPart2_l802 = (outPixelAddr_value % 3'b100);
  assign CICC1851_when_SuperResolutionPart2_l560 = (2'b10 * bufferWAddr_value);
  assign CICC1851_when_SuperResolutionPart2_l560_1 = {1'd0, outPixelAddr_value};
  assign CICC1851_when_SuperResolutionPart2_l602 = (2'b10 * bufferWAddr_value);
  assign CICC1851_when_SuperResolutionPart2_l602_1 = (CICC1851_when_SuperResolutionPart2_l602_2 + {1'b0,outPixelAddr_value});
  assign CICC1851_when_SuperResolutionPart2_l602_3 = {1'b0,2'b10};
  assign CICC1851_when_SuperResolutionPart2_l602_2 = {10'd0, CICC1851_when_SuperResolutionPart2_l602_3};
  assign CICC1851_when_SuperResolutionPart2_l603 = (2'b10 * bufferWAddr_value);
  assign CICC1851_when_SuperResolutionPart2_l603_1 = {1'd0, outPixelAddr_value};
  assign CICC1851_when_SuperResolutionPart2_l605 = (2'b10 * bufferWAddr_value);
  assign CICC1851_when_SuperResolutionPart2_l605_1 = (CICC1851_when_SuperResolutionPart2_l605_2 + {1'b0,outPixelAddr_value});
  assign CICC1851_when_SuperResolutionPart2_l605_3 = {1'b0,2'b11};
  assign CICC1851_when_SuperResolutionPart2_l605_2 = {10'd0, CICC1851_when_SuperResolutionPart2_l605_3};
  assign CICC1851_when_SuperResolutionPart2_l606 = (2'b10 * bufferWAddr_value);
  assign CICC1851_when_SuperResolutionPart2_l606_1 = (CICC1851_when_SuperResolutionPart2_l606_2 + {1'b0,outPixelAddr_value});
  assign CICC1851_when_SuperResolutionPart2_l606_3 = {1'b0,1'b1};
  assign CICC1851_when_SuperResolutionPart2_l606_2 = {11'd0, CICC1851_when_SuperResolutionPart2_l606_3};
  assign CICC1851_when_SuperResolutionPart2_l609 = (outPixelAddr_value % 2'b10);
  assign CICC1851_mainAddrOne_1 = (CICC1851_mainAddrOne_2 / 2'b10);
  assign CICC1851_mainAddrOne_2 = (outPixelAddr_value - 12'h002);
  assign CICC1851_mainAddrTwo_1 = (CICC1851_mainAddrTwo_2 / 2'b10);
  assign CICC1851_mainAddrTwo_2 = (outPixelAddr_value - 12'h002);
  assign CICC1851_when_SuperResolutionPart2_l667 = (CICC1851_when_SuperResolutionPart2_l667_1 - 13'h0002);
  assign CICC1851_when_SuperResolutionPart2_l667_1 = (2'b10 * bufferWAddr_value);
  assign CICC1851_when_SuperResolutionPart2_l667_2 = (CICC1851_when_SuperResolutionPart2_l667_3 + {1'b0,outPixelAddr_value});
  assign CICC1851_when_SuperResolutionPart2_l667_4 = {1'b0,1'b1};
  assign CICC1851_when_SuperResolutionPart2_l667_3 = {11'd0, CICC1851_when_SuperResolutionPart2_l667_4};
  assign CICC1851_when_SuperResolutionPart2_l668 = (2'b10 * bufferWAddr_value);
  assign CICC1851_when_SuperResolutionPart2_l668_1 = (CICC1851_when_SuperResolutionPart2_l668_2 + {1'b0,outPixelAddr_value});
  assign CICC1851_when_SuperResolutionPart2_l668_3 = {1'b0,1'b1};
  assign CICC1851_when_SuperResolutionPart2_l668_2 = {11'd0, CICC1851_when_SuperResolutionPart2_l668_3};
  assign CICC1851_mainAddrOne_3 = (CICC1851_mainAddrOne_4 / 2'b10);
  assign CICC1851_mainAddrOne_4 = (outPixelAddr_value - 12'h002);
  assign CICC1851_mainAddrTwo_3 = (CICC1851_mainAddrTwo_4 / 2'b10);
  assign CICC1851_mainAddrTwo_4 = (outPixelAddr_value - 12'h002);
  assign CICC1851_controls_onceMode = 2'b10;
  assign CICC1851_controls_onceMode_1 = 2'b11;
  assign CICC1851_mainAddrOne_5 = (CICC1851_mainAddrOne_6 / 2'b10);
  assign CICC1851_mainAddrOne_6 = (outPixelAddr_value - 12'h003);
  assign CICC1851_counterAddrOne_1 = (CICC1851_counterAddrOne_2 / 2'b10);
  assign CICC1851_counterAddrOne_2 = (outPixelAddr_value - 12'h003);
  assign CICC1851_counterAddrOne_3 = (CICC1851_counterAddrOne_4 / 2'b10);
  assign CICC1851_counterAddrOne_4 = (12'h001 + outPixelAddr_value);
  assign CICC1851_controls_onceMode_2 = 1'b1;
  assign CICC1851_mainAddrTwo_5 = (CICC1851_mainAddrTwo_6 / 2'b10);
  assign CICC1851_mainAddrTwo_6 = (outPixelAddr_value - 12'h003);
  assign CICC1851_counterAddrTwo_1 = (CICC1851_counterAddrTwo_2 / 2'b10);
  assign CICC1851_counterAddrTwo_2 = (outPixelAddr_value - 12'h003);
  assign CICC1851_counterAddrTwo_3 = (CICC1851_counterAddrTwo_4 / 2'b10);
  assign CICC1851_counterAddrTwo_4 = (12'h001 + outPixelAddr_value);
  assign CICC1851_mainAddrOne_7 = (CICC1851_mainAddrOne_8 / 2'b10);
  assign CICC1851_mainAddrOne_8 = (outPixelAddr_value - 12'h003);
  assign CICC1851_mainAddrOne_9 = (CICC1851_mainAddrOne_10 / 2'b10);
  assign CICC1851_mainAddrOne_10 = (outPixelAddr_value - 12'h003);
  assign CICC1851_counterAddrOne_5 = (CICC1851_counterAddrOne_6 / 2'b10);
  assign CICC1851_counterAddrOne_6 = (CICC1851_counterAddrOne_7 + {1'b0,outPixelAddr_value});
  assign CICC1851_counterAddrOne_8 = {1'b0,1'b1};
  assign CICC1851_counterAddrOne_7 = {11'd0, CICC1851_counterAddrOne_8};
  assign CICC1851_controls_twiceMode = 2'b10;
  assign CICC1851_mainAddrTwo_7 = (CICC1851_mainAddrTwo_8 / 2'b10);
  assign CICC1851_mainAddrTwo_8 = (outPixelAddr_value - 12'h003);
  assign CICC1851_controls_twiceMode_1 = 2'b11;
  assign CICC1851_mainAddrTwo_9 = (CICC1851_mainAddrTwo_10 / 2'b10);
  assign CICC1851_mainAddrTwo_10 = (outPixelAddr_value - 12'h003);
  assign CICC1851_counterAddrTwo_5 = (CICC1851_counterAddrTwo_6 / 2'b10);
  assign CICC1851_counterAddrTwo_6 = (CICC1851_counterAddrTwo_7 + {1'b0,outPixelAddr_value});
  assign CICC1851_counterAddrTwo_8 = {1'b0,1'b1};
  assign CICC1851_counterAddrTwo_7 = {11'd0, CICC1851_counterAddrTwo_8};
  assign CICC1851_mainAddrOne_11 = (CICC1851_mainAddrOne_12 / 2'b10);
  assign CICC1851_mainAddrOne_12 = (outPixelAddr_value - 12'h003);
  assign CICC1851_counterAddrTwo_9 = (CICC1851_counterAddrTwo_10 / 2'b10);
  assign CICC1851_counterAddrTwo_10 = (outPixelAddr_value - 12'h003);
  assign CICC1851_mainAddrTwo_11 = (CICC1851_mainAddrTwo_12 / 2'b10);
  assign CICC1851_mainAddrTwo_12 = (outPixelAddr_value - 12'h003);
  assign CICC1851_counterAddrOne_9 = (CICC1851_counterAddrOne_10 / 2'b10);
  assign CICC1851_counterAddrOne_10 = (outPixelAddr_value - 12'h003);
  assign CICC1851_mainAddrTwo_13 = (CICC1851_mainAddrTwo_14 / 2'b10);
  assign CICC1851_mainAddrTwo_14 = ({1'b0,outPixelAddr_value} + CICC1851_mainAddrTwo_15);
  assign CICC1851_mainAddrTwo_16 = {1'b0,1'b1};
  assign CICC1851_mainAddrTwo_15 = {11'd0, CICC1851_mainAddrTwo_16};
  assign CICC1851_counterAddrOne_11 = (CICC1851_counterAddrOne_12 / 2'b10);
  assign CICC1851_counterAddrOne_12 = ({1'b0,outPixelAddr_value} + CICC1851_counterAddrOne_13);
  assign CICC1851_counterAddrOne_14 = {1'b0,1'b1};
  assign CICC1851_counterAddrOne_13 = {11'd0, CICC1851_counterAddrOne_14};
  assign CICC1851_controls_twiceMode_2 = 1'b1;
  assign CICC1851_mainAddrTwo_17 = (CICC1851_mainAddrTwo_18 / 2'b10);
  assign CICC1851_mainAddrTwo_18 = (outPixelAddr_value - 12'h003);
  assign CICC1851_counterAddrOne_15 = (CICC1851_counterAddrOne_16 / 2'b10);
  assign CICC1851_counterAddrOne_16 = (outPixelAddr_value - 12'h003);
  assign CICC1851_mainAddrOne_13 = (CICC1851_mainAddrOne_14 / 2'b10);
  assign CICC1851_mainAddrOne_14 = (outPixelAddr_value - 12'h003);
  assign CICC1851_counterAddrTwo_11 = (CICC1851_counterAddrTwo_12 / 2'b10);
  assign CICC1851_counterAddrTwo_12 = (outPixelAddr_value - 12'h003);
  assign CICC1851_mainAddrOne_15 = (CICC1851_mainAddrOne_16 / 2'b10);
  assign CICC1851_mainAddrOne_16 = ({1'b0,outPixelAddr_value} + CICC1851_mainAddrOne_17);
  assign CICC1851_mainAddrOne_18 = {1'b0,1'b1};
  assign CICC1851_mainAddrOne_17 = {11'd0, CICC1851_mainAddrOne_18};
  assign CICC1851_counterAddrTwo_13 = (CICC1851_counterAddrTwo_14 / 2'b10);
  assign CICC1851_counterAddrTwo_14 = ({1'b0,outPixelAddr_value} + CICC1851_counterAddrTwo_15);
  assign CICC1851_counterAddrTwo_16 = {1'b0,1'b1};
  assign CICC1851_counterAddrTwo_15 = {11'd0, CICC1851_counterAddrTwo_16};
  assign CICC1851_lineBufferOne_port = passPixels_payload_pixel;
  assign CICC1851_lineBufferOne_port_1 = (passPixels_fire_6 && (bufferSwitch == 2'b00));
  assign CICC1851_lineBufferTwo_port = passPixels_payload_pixel;
  assign CICC1851_lineBufferTwo_port_1 = (passPixels_fire_8 && (bufferSwitch == 2'b10));
  assign CICC1851_lineBufferOdd_port = passPixels_payload_pixel;
  assign CICC1851_lineBufferOdd_port_1 = (passPixels_fire_7 && (bufferSwitch == 2'b01));
  always @(posedge clk) begin
    if(CICC1851_lineBufferOne_port_1) begin
      lineBufferOne[bufferWAddr_value] <= CICC1851_lineBufferOne_port;
    end
  end

  always @(posedge clk) begin
    if(mainAddrOneStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferOne_port1 <= lineBufferOne[mainAddrOneStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(counterAddrOneStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferOne_port2 <= lineBufferOne[counterAddrOneStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(CICC1851_lineBufferTwo_port_1) begin
      lineBufferTwo[bufferWAddr_value] <= CICC1851_lineBufferTwo_port;
    end
  end

  always @(posedge clk) begin
    if(mainAddrTwoStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferTwo_port1 <= lineBufferTwo[mainAddrTwoStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(counterAddrTwoStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferTwo_port2 <= lineBufferTwo[counterAddrTwoStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(CICC1851_lineBufferOdd_port_1) begin
      lineBufferOdd[bufferWAddr_value] <= CICC1851_lineBufferOdd_port;
    end
  end

  always @(posedge clk) begin
    if(oddAddrStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferOdd_port1 <= lineBufferOdd[oddAddrStream_s2mPipe_m2sPipe_payload];
    end
  end

  StreamFork_2 diffStage_controlPipe_fork (
    .io_input_valid                      (diffStage_controlPipe_valid                                     ), //i
    .io_input_ready                      (diffStage_controlPipe_fork_io_input_ready                       ), //o
    .io_input_payload_frameStart         (diffStage_controlPipe_payload_frameStart                        ), //i
    .io_input_payload_rowEnd             (diffStage_controlPipe_payload_rowEnd                            ), //i
    .io_input_payload_passMode           (diffStage_controlPipe_payload_passMode                          ), //i
    .io_input_payload_passValid          (diffStage_controlPipe_payload_passValid                         ), //i
    .io_input_payload_onceMode           (diffStage_controlPipe_payload_onceMode[2:0]                     ), //i
    .io_input_payload_onceValid          (diffStage_controlPipe_payload_onceValid                         ), //i
    .io_input_payload_mainCompare        (diffStage_controlPipe_payload_mainCompare                       ), //i
    .io_input_payload_counterCompare     (diffStage_controlPipe_payload_counterCompare                    ), //i
    .io_input_payload_mainDiff           (diffStage_controlPipe_payload_mainDiff[7:0]                     ), //i
    .io_input_payload_counterDiff        (diffStage_controlPipe_payload_counterDiff[7:0]                  ), //i
    .io_input_payload_twiceCompValid     (diffStage_controlPipe_payload_twiceCompValid                    ), //i
    .io_input_payload_twiceMode          (diffStage_controlPipe_payload_twiceMode[2:0]                    ), //i
    .io_input_payload_inpValidFlag       (diffStage_controlPipe_payload_inpValidFlag                      ), //i
    .io_input_payload_oddValid           (diffStage_controlPipe_payload_oddValid                          ), //i
    .io_outputs_0_valid                  (diffStage_controlPipe_fork_io_outputs_0_valid                   ), //o
    .io_outputs_0_ready                  (diffStage_controlPipe_fork_io_outputs_0_translated_ready        ), //i
    .io_outputs_0_payload_frameStart     (diffStage_controlPipe_fork_io_outputs_0_payload_frameStart      ), //o
    .io_outputs_0_payload_rowEnd         (diffStage_controlPipe_fork_io_outputs_0_payload_rowEnd          ), //o
    .io_outputs_0_payload_passMode       (diffStage_controlPipe_fork_io_outputs_0_payload_passMode        ), //o
    .io_outputs_0_payload_passValid      (diffStage_controlPipe_fork_io_outputs_0_payload_passValid       ), //o
    .io_outputs_0_payload_onceMode       (diffStage_controlPipe_fork_io_outputs_0_payload_onceMode[2:0]   ), //o
    .io_outputs_0_payload_onceValid      (diffStage_controlPipe_fork_io_outputs_0_payload_onceValid       ), //o
    .io_outputs_0_payload_mainCompare    (diffStage_controlPipe_fork_io_outputs_0_payload_mainCompare     ), //o
    .io_outputs_0_payload_counterCompare (diffStage_controlPipe_fork_io_outputs_0_payload_counterCompare  ), //o
    .io_outputs_0_payload_mainDiff       (diffStage_controlPipe_fork_io_outputs_0_payload_mainDiff[7:0]   ), //o
    .io_outputs_0_payload_counterDiff    (diffStage_controlPipe_fork_io_outputs_0_payload_counterDiff[7:0]), //o
    .io_outputs_0_payload_twiceCompValid (diffStage_controlPipe_fork_io_outputs_0_payload_twiceCompValid  ), //o
    .io_outputs_0_payload_twiceMode      (diffStage_controlPipe_fork_io_outputs_0_payload_twiceMode[2:0]  ), //o
    .io_outputs_0_payload_inpValidFlag   (diffStage_controlPipe_fork_io_outputs_0_payload_inpValidFlag    ), //o
    .io_outputs_0_payload_oddValid       (diffStage_controlPipe_fork_io_outputs_0_payload_oddValid        ), //o
    .io_outputs_1_valid                  (diffStage_controlPipe_fork_io_outputs_1_valid                   ), //o
    .io_outputs_1_ready                  (resultStage_pixelStream_ready                                   ), //i
    .io_outputs_1_payload_frameStart     (diffStage_controlPipe_fork_io_outputs_1_payload_frameStart      ), //o
    .io_outputs_1_payload_rowEnd         (diffStage_controlPipe_fork_io_outputs_1_payload_rowEnd          ), //o
    .io_outputs_1_payload_passMode       (diffStage_controlPipe_fork_io_outputs_1_payload_passMode        ), //o
    .io_outputs_1_payload_passValid      (diffStage_controlPipe_fork_io_outputs_1_payload_passValid       ), //o
    .io_outputs_1_payload_onceMode       (diffStage_controlPipe_fork_io_outputs_1_payload_onceMode[2:0]   ), //o
    .io_outputs_1_payload_onceValid      (diffStage_controlPipe_fork_io_outputs_1_payload_onceValid       ), //o
    .io_outputs_1_payload_mainCompare    (diffStage_controlPipe_fork_io_outputs_1_payload_mainCompare     ), //o
    .io_outputs_1_payload_counterCompare (diffStage_controlPipe_fork_io_outputs_1_payload_counterCompare  ), //o
    .io_outputs_1_payload_mainDiff       (diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff[7:0]   ), //o
    .io_outputs_1_payload_counterDiff    (diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff[7:0]), //o
    .io_outputs_1_payload_twiceCompValid (diffStage_controlPipe_fork_io_outputs_1_payload_twiceCompValid  ), //o
    .io_outputs_1_payload_twiceMode      (diffStage_controlPipe_fork_io_outputs_1_payload_twiceMode[2:0]  ), //o
    .io_outputs_1_payload_inpValidFlag   (diffStage_controlPipe_fork_io_outputs_1_payload_inpValidFlag    ), //o
    .io_outputs_1_payload_oddValid       (diffStage_controlPipe_fork_io_outputs_1_payload_oddValid        )  //o
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_7_BOOT : controlStateMachine_stateReg_string = "BOOT ";
      controlStateMachine_enumDef_7_HOLD : controlStateMachine_stateReg_string = "HOLD ";
      controlStateMachine_enumDef_7_PASS : controlStateMachine_stateReg_string = "PASS ";
      controlStateMachine_enumDef_7_ONCE : controlStateMachine_stateReg_string = "ONCE ";
      controlStateMachine_enumDef_7_TWICE : controlStateMachine_stateReg_string = "TWICE";
      default : controlStateMachine_stateReg_string = "?????";
    endcase
  end
  always @(*) begin
    case(controlStateMachine_stateNext)
      controlStateMachine_enumDef_7_BOOT : controlStateMachine_stateNext_string = "BOOT ";
      controlStateMachine_enumDef_7_HOLD : controlStateMachine_stateNext_string = "HOLD ";
      controlStateMachine_enumDef_7_PASS : controlStateMachine_stateNext_string = "PASS ";
      controlStateMachine_enumDef_7_ONCE : controlStateMachine_stateNext_string = "ONCE ";
      controlStateMachine_enumDef_7_TWICE : controlStateMachine_stateNext_string = "TWICE";
      default : controlStateMachine_stateNext_string = "?????";
    endcase
  end
  `endif

  always @(*) begin
    pixelsIn_ready = 1'b0;
    pixelsIn_ready = (! pixelsIn_rValid);
  end

  always @(*) begin
    pixelsOut_valid = 1'b0;
    pixelsOut_valid = pixelsStream_s2mPipe_m2sPipe_valid;
  end

  always @(*) begin
    pixelsOut_payload_pixel = 8'h0;
    pixelsOut_payload_pixel = pixelsStream_s2mPipe_m2sPipe_payload_pixel;
  end

  always @(*) begin
    pixelsOut_payload_frameStart = 1'b0;
    pixelsOut_payload_frameStart = pixelsStream_s2mPipe_m2sPipe_payload_frameStart;
  end

  always @(*) begin
    pixelsOut_payload_rowEnd = 1'b0;
    pixelsOut_payload_rowEnd = pixelsStream_s2mPipe_m2sPipe_payload_rowEnd;
  end

  always @(*) begin
    pixelsOut_payload_inpValid = 1'b0;
    pixelsOut_payload_inpValid = pixelsStream_s2mPipe_m2sPipe_payload_inpValid;
  end

  always @(*) begin
    startOut = 1'b0;
    startOut = slaveStart;
  end

  always @(*) begin
    inpTwoDoneOut = 1'b0;
    inpTwoDoneOut = inpTwoDone;
  end

  assign when_SuperResolutionPart2_l40 = (inpThreeDoneIn || (startIn && (! startIn_regNext)));
  assign when_SuperResolutionPart2_l43 = (! startIn);
  assign when_SuperResolutionPart2_l46 = (startIn && (! readDone));
  assign when_SuperResolutionPart2_l46_1 = (! startIn);
  assign pixelsIn_fire = (pixelsIn_valid && pixelsIn_ready);
  assign when_SuperResolutionPart2_l49 = ((! inpThreeDoneIn) && pixelsIn_fire);
  assign when_SuperResolutionPart2_l49_1 = (inpThreeDoneIn || (! startIn));
  assign when_SuperResolutionPart2_l64 = (! startIn);
  assign when_SuperResolutionPart2_l67 = (! startIn);
  always @(*) begin
    bufferRowCount_willIncrement = 1'b0;
    if(when_SuperResolutionPart2_l185) begin
      if(!bufferReachFinalRow) begin
        bufferRowCount_willIncrement = 1'b1;
      end
    end
  end

  always @(*) begin
    bufferRowCount_willClear = 1'b0;
    if(when_SuperResolutionPart2_l185) begin
      if(bufferReachFinalRow) begin
        bufferRowCount_willClear = 1'b1;
      end
    end
  end

  assign bufferRowCount_willOverflowIfInc = (bufferRowCount_value == 11'h438);
  assign bufferRowCount_willOverflow = (bufferRowCount_willOverflowIfInc && bufferRowCount_willIncrement);
  always @(*) begin
    if(bufferRowCount_willOverflow) begin
      bufferRowCount_valueNext = 11'h0;
    end else begin
      bufferRowCount_valueNext = (bufferRowCount_value + CICC1851_bufferRowCount_valueNext);
    end
    if(bufferRowCount_willClear) begin
      bufferRowCount_valueNext = 11'h0;
    end
  end

  assign when_SuperResolutionPart2_l76 = ((startIn && (! holdBuffer)) && (! writeDone));
  assign when_SuperResolutionPart2_l76_1 = (((! startIn) || holdBuffer) || writeDone);
  assign when_SuperResolutionPart2_l82 = (! startRead);
  always @(*) begin
    bufferWAddr_willIncrement = 1'b0;
    if(passPixels_fire_9) begin
      if(!passPixels_payload_rowEnd) begin
        bufferWAddr_willIncrement = 1'b1;
      end
    end
  end

  always @(*) begin
    bufferWAddr_willClear = 1'b0;
    if(passPixels_fire_9) begin
      if(passPixels_payload_rowEnd) begin
        bufferWAddr_willClear = 1'b1;
      end
    end
  end

  assign bufferWAddr_willOverflowIfInc = (bufferWAddr_value == 11'h77f);
  assign bufferWAddr_willOverflow = (bufferWAddr_willOverflowIfInc && bufferWAddr_willIncrement);
  always @(*) begin
    if(bufferWAddr_willOverflow) begin
      bufferWAddr_valueNext = 11'h0;
    end else begin
      bufferWAddr_valueNext = (bufferWAddr_value + CICC1851_bufferWAddr_valueNext);
    end
    if(bufferWAddr_willClear) begin
      bufferWAddr_valueNext = 11'h0;
    end
  end

  always @(*) begin
    outPixelAddr_willIncrement = 1'b0;
    if(when_SuperResolutionPart2_l761) begin
      if(controlStream_fire_7) begin
        if(!outReachRowEnd) begin
          outPixelAddr_willIncrement = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    outPixelAddr_willClear = 1'b0;
    if(when_SuperResolutionPart2_l761) begin
      if(controlStream_fire_7) begin
        if(outReachRowEnd) begin
          outPixelAddr_willClear = 1'b1;
        end
      end
    end
  end

  assign outPixelAddr_willOverflowIfInc = (outPixelAddr_value == 12'heff);
  assign outPixelAddr_willOverflow = (outPixelAddr_willOverflowIfInc && outPixelAddr_willIncrement);
  always @(*) begin
    if(outPixelAddr_willOverflow) begin
      outPixelAddr_valueNext = 12'h0;
    end else begin
      outPixelAddr_valueNext = (outPixelAddr_value + CICC1851_outPixelAddr_valueNext);
    end
    if(outPixelAddr_willClear) begin
      outPixelAddr_valueNext = 12'h0;
    end
  end

  always @(*) begin
    outRowCount_willIncrement = 1'b0;
    if(when_SuperResolutionPart2_l761) begin
      if(when_SuperResolutionPart2_l766) begin
        if(!outReachFinalRow) begin
          outRowCount_willIncrement = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    outRowCount_willClear = 1'b0;
    if(when_SuperResolutionPart2_l761) begin
      if(when_SuperResolutionPart2_l766) begin
        if(outReachFinalRow) begin
          outRowCount_willClear = 1'b1;
        end
      end
    end
  end

  assign outRowCount_willOverflowIfInc = (outRowCount_value == 12'h870);
  assign outRowCount_willOverflow = (outRowCount_willOverflowIfInc && outRowCount_willIncrement);
  always @(*) begin
    if(outRowCount_willOverflow) begin
      outRowCount_valueNext = 12'h0;
    end else begin
      outRowCount_valueNext = (outRowCount_value + CICC1851_outRowCount_valueNext);
    end
    if(outRowCount_willClear) begin
      outRowCount_valueNext = 12'h0;
    end
  end

  always @(*) begin
    alreadySendRow_willIncrement = 1'b0;
    if(pixelsOut_fire_2) begin
      if(alreadyReachRowEnd) begin
        if(!alreadyReachFinalRow) begin
          alreadySendRow_willIncrement = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    alreadySendRow_willClear = 1'b0;
    if(pixelsOut_fire_2) begin
      if(alreadyReachRowEnd) begin
        if(alreadyReachFinalRow) begin
          alreadySendRow_willClear = 1'b1;
        end
      end
    end
  end

  assign alreadySendRow_willOverflowIfInc = (alreadySendRow_value == 12'h870);
  assign alreadySendRow_willOverflow = (alreadySendRow_willOverflowIfInc && alreadySendRow_willIncrement);
  always @(*) begin
    if(alreadySendRow_willOverflow) begin
      alreadySendRow_valueNext = 12'h0;
    end else begin
      alreadySendRow_valueNext = (alreadySendRow_value + CICC1851_alreadySendRow_valueNext);
    end
    if(alreadySendRow_willClear) begin
      alreadySendRow_valueNext = 12'h0;
    end
  end

  always @(*) begin
    alreadySendCountInRow_willIncrement = 1'b0;
    if(pixelsOut_fire_2) begin
      if(!alreadyReachRowEnd) begin
        alreadySendCountInRow_willIncrement = 1'b1;
      end
    end
  end

  always @(*) begin
    alreadySendCountInRow_willClear = 1'b0;
    if(pixelsOut_fire_2) begin
      if(alreadyReachRowEnd) begin
        alreadySendCountInRow_willClear = 1'b1;
      end
    end
  end

  assign alreadySendCountInRow_willOverflowIfInc = (alreadySendCountInRow_value == 12'heff);
  assign alreadySendCountInRow_willOverflow = (alreadySendCountInRow_willOverflowIfInc && alreadySendCountInRow_willIncrement);
  always @(*) begin
    if(alreadySendCountInRow_willOverflow) begin
      alreadySendCountInRow_valueNext = 12'h0;
    end else begin
      alreadySendCountInRow_valueNext = (alreadySendCountInRow_value + CICC1851_alreadySendCountInRow_valueNext);
    end
    if(alreadySendCountInRow_willClear) begin
      alreadySendCountInRow_valueNext = 12'h0;
    end
  end

  assign when_SuperResolutionPart2_l106 = (((! startIn) && startIn_regNext_1) || inpTwoDone);
  assign when_SuperResolutionPart2_l108 = (((! startIn) && startIn_regNext_2) || inpTwoDone);
  assign when_SuperResolutionPart2_l109 = (((! startIn) && startIn_regNext_3) || inpTwoDone);
  assign when_SuperResolutionPart2_l110 = (((! startIn) && startIn_regNext_4) || inpTwoDone);
  assign when_SuperResolutionPart2_l111 = (((! startIn) && startIn_regNext_5) || inpTwoDone);
  assign when_SuperResolutionPart2_l113 = (((! startIn) && startIn_regNext_6) || inpTwoDone);
  assign when_SuperResolutionPart2_l114 = (((! startIn) && startIn_regNext_7) || inpTwoDone);
  assign when_SuperResolutionPart2_l115 = (((! startIn) && startIn_regNext_8) || inpTwoDone);
  assign when_SuperResolutionPart2_l116 = (((! startIn) && startIn_regNext_9) || inpTwoDone);
  assign when_SuperResolutionPart2_l120 = (((! startIn) && startIn_regNext_10) || inpTwoDone);
  assign when_SuperResolutionPart2_l121 = (((! startIn) && startIn_regNext_11) || inpTwoDone);
  assign when_SuperResolutionPart2_l122 = (((! startIn) && startIn_regNext_12) || inpTwoDone);
  assign when_SuperResolutionPart2_l123 = (((! startIn) && startIn_regNext_13) || inpTwoDone);
  assign when_SuperResolutionPart2_l124 = (((! startIn) && startIn_regNext_14) || inpTwoDone);
  assign when_SuperResolutionPart2_l125 = (((! startIn) && startIn_regNext_15) || inpTwoDone);
  assign when_SuperResolutionPart2_l126 = (((! startIn) && startIn_regNext_16) || inpTwoDone);
  assign when_SuperResolutionPart2_l134 = (! startRead);
  always @(*) begin
    mainAddrOne = CICC1851_mainAddrOne[10:0];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_7_HOLD : begin
      end
      controlStateMachine_enumDef_7_PASS : begin
        if(!twoInFourOutRow) begin
          if(oneInFourOutRow) begin
            if(nextRowBuffer) begin
              if(twoInFourOutPixelAddr) begin
                mainAddrOne = CICC1851_mainAddrOne_1[10:0];
              end
            end
          end
        end
      end
      controlStateMachine_enumDef_7_ONCE : begin
        if(threeInFourOutRow) begin
          if(twoInFourOutPixelAddr) begin
            mainAddrOne = CICC1851_mainAddrOne_3[10:0];
          end
        end else begin
          if(nextRowBuffer) begin
            mainAddrOne = CICC1851_mainAddrOne_5[10:0];
          end
        end
      end
      controlStateMachine_enumDef_7_TWICE : begin
        if(outReachFinalRow) begin
          if(nextRowBuffer) begin
            if(outReachRowEnd) begin
              mainAddrOne = CICC1851_mainAddrOne_7[10:0];
            end else begin
              mainAddrOne = CICC1851_mainAddrOne_9[10:0];
            end
          end
        end else begin
          if(nextRowBuffer) begin
            mainAddrOne = CICC1851_mainAddrOne_11[10:0];
          end else begin
            if(outReachRowEnd) begin
              mainAddrOne = CICC1851_mainAddrOne_13[10:0];
            end else begin
              mainAddrOne = CICC1851_mainAddrOne_15[10:0];
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    counterAddrOne = CICC1851_counterAddrOne[10:0];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_7_HOLD : begin
      end
      controlStateMachine_enumDef_7_PASS : begin
      end
      controlStateMachine_enumDef_7_ONCE : begin
        if(!threeInFourOutRow) begin
          if(nextRowBuffer) begin
            if(outReachRowEnd) begin
              counterAddrOne = CICC1851_counterAddrOne_1[10:0];
            end else begin
              counterAddrOne = CICC1851_counterAddrOne_3[10:0];
            end
          end
        end
      end
      controlStateMachine_enumDef_7_TWICE : begin
        if(outReachFinalRow) begin
          if(nextRowBuffer) begin
            if(!outReachRowEnd) begin
              counterAddrOne = CICC1851_counterAddrOne_5[10:0];
            end
          end
        end else begin
          if(nextRowBuffer) begin
            if(outReachRowEnd) begin
              counterAddrOne = CICC1851_counterAddrOne_9[10:0];
            end else begin
              counterAddrOne = CICC1851_counterAddrOne_11[10:0];
            end
          end else begin
            counterAddrOne = CICC1851_counterAddrOne_15[10:0];
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    mainAddrTwo = CICC1851_mainAddrTwo[10:0];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_7_HOLD : begin
      end
      controlStateMachine_enumDef_7_PASS : begin
        if(!twoInFourOutRow) begin
          if(oneInFourOutRow) begin
            if(!nextRowBuffer) begin
              if(twoInFourOutPixelAddr) begin
                mainAddrTwo = CICC1851_mainAddrTwo_1[10:0];
              end
            end
          end
        end
      end
      controlStateMachine_enumDef_7_ONCE : begin
        if(threeInFourOutRow) begin
          if(twoInFourOutPixelAddr) begin
            mainAddrTwo = CICC1851_mainAddrTwo_3[10:0];
          end
        end else begin
          if(!nextRowBuffer) begin
            mainAddrTwo = CICC1851_mainAddrTwo_5[10:0];
          end
        end
      end
      controlStateMachine_enumDef_7_TWICE : begin
        if(outReachFinalRow) begin
          if(!nextRowBuffer) begin
            if(outReachRowEnd) begin
              mainAddrTwo = CICC1851_mainAddrTwo_7[10:0];
            end else begin
              mainAddrTwo = CICC1851_mainAddrTwo_9[10:0];
            end
          end
        end else begin
          if(nextRowBuffer) begin
            if(outReachRowEnd) begin
              mainAddrTwo = CICC1851_mainAddrTwo_11[10:0];
            end else begin
              mainAddrTwo = CICC1851_mainAddrTwo_13[10:0];
            end
          end else begin
            mainAddrTwo = CICC1851_mainAddrTwo_17[10:0];
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    counterAddrTwo = CICC1851_counterAddrTwo[10:0];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_7_HOLD : begin
      end
      controlStateMachine_enumDef_7_PASS : begin
      end
      controlStateMachine_enumDef_7_ONCE : begin
        if(!threeInFourOutRow) begin
          if(!nextRowBuffer) begin
            if(outReachRowEnd) begin
              counterAddrTwo = CICC1851_counterAddrTwo_1[10:0];
            end else begin
              counterAddrTwo = CICC1851_counterAddrTwo_3[10:0];
            end
          end
        end
      end
      controlStateMachine_enumDef_7_TWICE : begin
        if(outReachFinalRow) begin
          if(!nextRowBuffer) begin
            if(!outReachRowEnd) begin
              counterAddrTwo = CICC1851_counterAddrTwo_5[10:0];
            end
          end
        end else begin
          if(nextRowBuffer) begin
            counterAddrTwo = CICC1851_counterAddrTwo_9[10:0];
          end else begin
            if(outReachRowEnd) begin
              counterAddrTwo = CICC1851_counterAddrTwo_11[10:0];
            end else begin
              counterAddrTwo = CICC1851_counterAddrTwo_13[10:0];
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign oddAddr = CICC1851_oddAddr[10:0];
  assign validStream_valid = 1'b1;
  assign CICC1851_controls_frameStart = 32'h0;
  always @(*) begin
    controls_frameStart = CICC1851_controls_frameStart[0];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_7_HOLD : begin
      end
      controlStateMachine_enumDef_7_PASS : begin
        if(frameStart) begin
          controls_frameStart = 1'b1;
        end
      end
      controlStateMachine_enumDef_7_ONCE : begin
      end
      controlStateMachine_enumDef_7_TWICE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_rowEnd = CICC1851_controls_frameStart[1];
    if(when_SuperResolutionPart2_l761) begin
      if(outReachRowEnd) begin
        controls_rowEnd = 1'b1;
      end
    end
  end

  always @(*) begin
    controls_passMode = CICC1851_controls_frameStart[2];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_7_HOLD : begin
      end
      controlStateMachine_enumDef_7_PASS : begin
        if(twoInFourOutRow) begin
          if(!when_SuperResolutionPart2_l609) begin
            if(nextRowBuffer) begin
              controls_passMode = 1'b0;
            end else begin
              controls_passMode = 1'b1;
            end
          end
        end else begin
          if(oneInFourOutRow) begin
            if(nextRowBuffer) begin
              controls_passMode = 1'b0;
            end else begin
              controls_passMode = 1'b1;
            end
          end else begin
            if(nextRowBuffer) begin
              controls_passMode = 1'b0;
            end else begin
              controls_passMode = 1'b1;
            end
          end
        end
      end
      controlStateMachine_enumDef_7_ONCE : begin
      end
      controlStateMachine_enumDef_7_TWICE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_passValid = CICC1851_controls_frameStart[3];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_7_HOLD : begin
      end
      controlStateMachine_enumDef_7_PASS : begin
        if(twoInFourOutRow) begin
          if(!when_SuperResolutionPart2_l609) begin
            controls_passValid = 1'b1;
          end
        end else begin
          if(oneInFourOutRow) begin
            controls_passValid = 1'b1;
          end else begin
            controls_passValid = 1'b1;
          end
        end
      end
      controlStateMachine_enumDef_7_ONCE : begin
      end
      controlStateMachine_enumDef_7_TWICE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_onceMode = CICC1851_controls_frameStart[6 : 4];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_7_HOLD : begin
      end
      controlStateMachine_enumDef_7_PASS : begin
      end
      controlStateMachine_enumDef_7_ONCE : begin
        if(threeInFourOutRow) begin
          if(outReachFinalRow) begin
            if(nextRowBuffer) begin
              controls_onceMode = 3'b100;
            end else begin
              controls_onceMode = 3'b101;
            end
          end else begin
            if(nextRowBuffer) begin
              controls_onceMode = {1'd0, CICC1851_controls_onceMode};
            end else begin
              controls_onceMode = {1'd0, CICC1851_controls_onceMode_1};
            end
          end
        end else begin
          if(nextRowBuffer) begin
            controls_onceMode = 3'b000;
          end else begin
            controls_onceMode = {2'd0, CICC1851_controls_onceMode_2};
          end
        end
      end
      controlStateMachine_enumDef_7_TWICE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_onceValid = CICC1851_controls_frameStart[7];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_7_HOLD : begin
      end
      controlStateMachine_enumDef_7_PASS : begin
      end
      controlStateMachine_enumDef_7_ONCE : begin
        controls_onceValid = 1'b1;
      end
      controlStateMachine_enumDef_7_TWICE : begin
      end
      default : begin
      end
    endcase
  end

  assign controls_mainCompare = CICC1851_controls_frameStart[8];
  assign controls_counterCompare = CICC1851_controls_frameStart[9];
  assign controls_mainDiff = CICC1851_controls_frameStart[17 : 10];
  assign controls_counterDiff = CICC1851_controls_frameStart[25 : 18];
  always @(*) begin
    controls_twiceCompValid = CICC1851_controls_frameStart[26];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_7_HOLD : begin
      end
      controlStateMachine_enumDef_7_PASS : begin
      end
      controlStateMachine_enumDef_7_ONCE : begin
      end
      controlStateMachine_enumDef_7_TWICE : begin
        controls_twiceCompValid = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_twiceMode = CICC1851_controls_frameStart[29 : 27];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_7_HOLD : begin
      end
      controlStateMachine_enumDef_7_PASS : begin
      end
      controlStateMachine_enumDef_7_ONCE : begin
      end
      controlStateMachine_enumDef_7_TWICE : begin
        if(outReachFinalRow) begin
          if(nextRowBuffer) begin
            if(outReachRowEnd) begin
              controls_twiceMode = 3'b100;
            end else begin
              controls_twiceMode = 3'b101;
            end
          end else begin
            if(outReachRowEnd) begin
              controls_twiceMode = {1'd0, CICC1851_controls_twiceMode};
            end else begin
              controls_twiceMode = {1'd0, CICC1851_controls_twiceMode_1};
            end
          end
        end else begin
          if(nextRowBuffer) begin
            controls_twiceMode = 3'b000;
          end else begin
            controls_twiceMode = {2'd0, CICC1851_controls_twiceMode_2};
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_inpValidFlag = CICC1851_controls_frameStart[30];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_7_HOLD : begin
        controls_inpValidFlag = 1'b1;
      end
      controlStateMachine_enumDef_7_PASS : begin
        controls_inpValidFlag = 1'b1;
      end
      controlStateMachine_enumDef_7_ONCE : begin
        controls_inpValidFlag = 1'b1;
      end
      controlStateMachine_enumDef_7_TWICE : begin
        controls_inpValidFlag = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_oddValid = CICC1851_controls_frameStart[31];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_7_HOLD : begin
      end
      controlStateMachine_enumDef_7_PASS : begin
        if(twoInFourOutRow) begin
          if(when_SuperResolutionPart2_l609) begin
            controls_oddValid = 1'b1;
          end
        end
      end
      controlStateMachine_enumDef_7_ONCE : begin
      end
      controlStateMachine_enumDef_7_TWICE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    validStream_ready = (controlStream_ready && startRead);
    validStream_ready = (mainAddrOneStream_ready && startRead);
    validStream_ready = (counterAddrOneStream_ready && startRead);
    validStream_ready = (mainAddrTwoStream_ready && startRead);
    validStream_ready = (counterAddrTwoStream_ready && startRead);
    validStream_ready = (oddAddrStream_ready && startRead);
  end

  assign controlStream_valid = (validStream_valid && startRead);
  assign controlStream_payload_frameStart = controls_frameStart;
  assign controlStream_payload_rowEnd = controls_rowEnd;
  assign controlStream_payload_passMode = controls_passMode;
  assign controlStream_payload_passValid = controls_passValid;
  assign controlStream_payload_onceMode = controls_onceMode;
  assign controlStream_payload_onceValid = controls_onceValid;
  assign controlStream_payload_mainCompare = controls_mainCompare;
  assign controlStream_payload_counterCompare = controls_counterCompare;
  assign controlStream_payload_mainDiff = controls_mainDiff;
  assign controlStream_payload_counterDiff = controls_counterDiff;
  assign controlStream_payload_twiceCompValid = controls_twiceCompValid;
  assign controlStream_payload_twiceMode = controls_twiceMode;
  assign controlStream_payload_inpValidFlag = controls_inpValidFlag;
  assign controlStream_payload_oddValid = controls_oddValid;
  assign mainAddrOneStream_valid = (validStream_valid && startRead);
  assign mainAddrOneStream_payload = mainAddrOne;
  assign counterAddrOneStream_valid = (validStream_valid && startRead);
  assign counterAddrOneStream_payload = counterAddrOne;
  assign mainAddrTwoStream_valid = (validStream_valid && startRead);
  assign mainAddrTwoStream_payload = mainAddrTwo;
  assign counterAddrTwoStream_valid = (validStream_valid && startRead);
  assign counterAddrTwoStream_payload = counterAddrTwo;
  assign oddAddrStream_valid = (validStream_valid && startRead);
  assign oddAddrStream_payload = oddAddr;
  assign pixelsIn_s2mPipe_valid = (pixelsIn_valid || pixelsIn_rValid);
  assign pixelsIn_s2mPipe_payload_pixel = (pixelsIn_rValid ? pixelsIn_rData_pixel : pixelsIn_payload_pixel);
  assign pixelsIn_s2mPipe_payload_frameStart = (pixelsIn_rValid ? pixelsIn_rData_frameStart : pixelsIn_payload_frameStart);
  assign pixelsIn_s2mPipe_payload_rowEnd = (pixelsIn_rValid ? pixelsIn_rData_rowEnd : pixelsIn_payload_rowEnd);
  always @(*) begin
    pixelsIn_s2mPipe_ready = pixelsIn_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368) begin
      pixelsIn_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368 = (! pixelsIn_s2mPipe_m2sPipe_valid);
  assign pixelsIn_s2mPipe_m2sPipe_valid = pixelsIn_s2mPipe_rValid;
  assign pixelsIn_s2mPipe_m2sPipe_payload_pixel = pixelsIn_s2mPipe_rData_pixel;
  assign pixelsIn_s2mPipe_m2sPipe_payload_frameStart = pixelsIn_s2mPipe_rData_frameStart;
  assign pixelsIn_s2mPipe_m2sPipe_payload_rowEnd = pixelsIn_s2mPipe_rData_rowEnd;
  assign passPixels_valid = (pixelsIn_s2mPipe_m2sPipe_valid && bufferEnable);
  assign pixelsIn_s2mPipe_m2sPipe_ready = (passPixels_ready && bufferEnable);
  assign passPixels_payload_pixel = pixelsIn_s2mPipe_m2sPipe_payload_pixel;
  assign passPixels_payload_frameStart = pixelsIn_s2mPipe_m2sPipe_payload_frameStart;
  assign passPixels_payload_rowEnd = pixelsIn_s2mPipe_m2sPipe_payload_rowEnd;
  assign passPixels_ready = 1'b1;
  assign passPixels_fire = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart2_l181 = ((CICC1851_when_SuperResolutionPart2_l181 == CICC1851_when_SuperResolutionPart2_l181_1) && passPixels_fire);
  assign passPixels_fire_1 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart2_l182 = (((CICC1851_when_SuperResolutionPart2_l182 == CICC1851_when_SuperResolutionPart2_l182_1) && bufferReachRowEnd) && passPixels_fire_1);
  assign passPixels_fire_2 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart2_l185 = (passPixels_payload_rowEnd && passPixels_fire_2);
  assign when_SuperResolutionPart2_l195 = (CICC1851_when_SuperResolutionPart2_l195 == 11'h0);
  assign passPixels_fire_3 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart2_l200 = (passPixels_payload_rowEnd && passPixels_fire_3);
  assign when_SuperResolutionPart2_l201 = ((bufferSwitch == 2'b10) || (bufferSwitch == 2'b00));
  assign passPixels_fire_4 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart2_l207 = (((bufferRowCount_value != 11'h0) && passPixels_payload_rowEnd) && passPixels_fire_4);
  assign when_SuperResolutionPart2_l208 = (bufferSwitch != 2'b01);
  assign when_SuperResolutionPart2_l212 = (bufferReachFinalRow && bufferReachRowEnd);
  assign controlStream_fire = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart2_l218 = (((CICC1851_when_SuperResolutionPart2_l218 == 12'h003) && controlStream_payload_rowEnd) && controlStream_fire);
  assign when_SuperResolutionPart2_l220 = 1'b1;
  assign passPixels_fire_5 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart2_l224 = (passPixels_payload_frameStart && passPixels_fire_5);
  assign pixelsOut_fire = (pixelsOut_valid && pixelsOut_ready);
  assign when_SuperResolutionPart2_l234 = ((CICC1851_when_SuperResolutionPart2_l234 == CICC1851_when_SuperResolutionPart2_l234_1) && pixelsOut_fire);
  assign pixelsOut_fire_1 = (pixelsOut_valid && pixelsOut_ready);
  assign when_SuperResolutionPart2_l235 = (((CICC1851_when_SuperResolutionPart2_l235 == CICC1851_when_SuperResolutionPart2_l235_1) && alreadyReachRowEnd) && pixelsOut_fire_1);
  assign pixelsOut_fire_2 = (pixelsOut_valid && pixelsOut_ready);
  assign pixelsOut_fire_3 = (pixelsOut_valid && pixelsOut_ready);
  assign when_SuperResolutionPart2_l246 = ((alreadyReachFinalRow && alreadyReachRowEnd) && pixelsOut_fire_3);
  assign passPixels_fire_6 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_7 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_8 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_9 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_10 = (passPixels_valid && passPixels_ready);
  assign controlStream_fire_1 = (controlStream_valid && controlStream_ready);
  assign pushing = (passPixels_fire_10 && (! controlStream_fire_1));
  assign passPixels_fire_11 = (passPixels_valid && passPixels_ready);
  assign controlStream_fire_2 = (controlStream_valid && controlStream_ready);
  assign poping = ((! passPixels_fire_11) && controlStream_fire_2);
  assign passPixels_fire_12 = (passPixels_valid && passPixels_ready);
  assign controlStream_fire_3 = (controlStream_valid && controlStream_ready);
  assign pushAndPoping = (passPixels_fire_12 && controlStream_fire_3);
  assign mainAddrOneStream_ready = (! mainAddrOneStream_rValid);
  assign mainAddrOneStream_s2mPipe_valid = (mainAddrOneStream_valid || mainAddrOneStream_rValid);
  assign mainAddrOneStream_s2mPipe_payload = (mainAddrOneStream_rValid ? mainAddrOneStream_rData : mainAddrOneStream_payload);
  always @(*) begin
    mainAddrOneStream_s2mPipe_ready = mainAddrOneStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_1) begin
      mainAddrOneStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_1 = (! mainAddrOneStream_s2mPipe_m2sPipe_valid);
  assign mainAddrOneStream_s2mPipe_m2sPipe_valid = mainAddrOneStream_s2mPipe_rValid;
  assign mainAddrOneStream_s2mPipe_m2sPipe_payload = mainAddrOneStream_s2mPipe_rData;
  assign mainAddrOneStream_s2mPipe_m2sPipe_ready = ((! CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready) || CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready = CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_mainOnePixelStream_payload = CICC1851_lineBufferOne_port1;
  assign CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_1 = readStage_mainOnePixelStream_ready;
    if(when_Stream_l368_2) begin
      CICC1851_1 = 1'b1;
    end
  end

  assign when_Stream_l368_2 = (! readStage_mainOnePixelStream_valid);
  assign readStage_mainOnePixelStream_valid = CICC1851_readStage_mainOnePixelStream_valid;
  assign readStage_mainOnePixelStream_payload = CICC1851_readStage_mainOnePixelStream_payload_2;
  assign counterAddrOneStream_ready = (! counterAddrOneStream_rValid);
  assign counterAddrOneStream_s2mPipe_valid = (counterAddrOneStream_valid || counterAddrOneStream_rValid);
  assign counterAddrOneStream_s2mPipe_payload = (counterAddrOneStream_rValid ? counterAddrOneStream_rData : counterAddrOneStream_payload);
  always @(*) begin
    counterAddrOneStream_s2mPipe_ready = counterAddrOneStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_3) begin
      counterAddrOneStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_3 = (! counterAddrOneStream_s2mPipe_m2sPipe_valid);
  assign counterAddrOneStream_s2mPipe_m2sPipe_valid = counterAddrOneStream_s2mPipe_rValid;
  assign counterAddrOneStream_s2mPipe_m2sPipe_payload = counterAddrOneStream_s2mPipe_rData;
  assign counterAddrOneStream_s2mPipe_m2sPipe_ready = ((! CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready) || CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready = CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_counterOnePixelStream_payload = CICC1851_lineBufferOne_port2;
  assign CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_2 = readStage_counterOnePixelStream_ready;
    if(when_Stream_l368_4) begin
      CICC1851_2 = 1'b1;
    end
  end

  assign when_Stream_l368_4 = (! readStage_counterOnePixelStream_valid);
  assign readStage_counterOnePixelStream_valid = CICC1851_readStage_counterOnePixelStream_valid;
  assign readStage_counterOnePixelStream_payload = CICC1851_readStage_counterOnePixelStream_payload_2;
  assign mainAddrTwoStream_ready = (! mainAddrTwoStream_rValid);
  assign mainAddrTwoStream_s2mPipe_valid = (mainAddrTwoStream_valid || mainAddrTwoStream_rValid);
  assign mainAddrTwoStream_s2mPipe_payload = (mainAddrTwoStream_rValid ? mainAddrTwoStream_rData : mainAddrTwoStream_payload);
  always @(*) begin
    mainAddrTwoStream_s2mPipe_ready = mainAddrTwoStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_5) begin
      mainAddrTwoStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_5 = (! mainAddrTwoStream_s2mPipe_m2sPipe_valid);
  assign mainAddrTwoStream_s2mPipe_m2sPipe_valid = mainAddrTwoStream_s2mPipe_rValid;
  assign mainAddrTwoStream_s2mPipe_m2sPipe_payload = mainAddrTwoStream_s2mPipe_rData;
  assign mainAddrTwoStream_s2mPipe_m2sPipe_ready = ((! CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready) || CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready = CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_mainTwoPixelStream_payload = CICC1851_lineBufferTwo_port1;
  assign CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_3 = readStage_mainTwoPixelStream_ready;
    if(when_Stream_l368_6) begin
      CICC1851_3 = 1'b1;
    end
  end

  assign when_Stream_l368_6 = (! readStage_mainTwoPixelStream_valid);
  assign readStage_mainTwoPixelStream_valid = CICC1851_readStage_mainTwoPixelStream_valid;
  assign readStage_mainTwoPixelStream_payload = CICC1851_readStage_mainTwoPixelStream_payload_2;
  assign counterAddrTwoStream_ready = (! counterAddrTwoStream_rValid);
  assign counterAddrTwoStream_s2mPipe_valid = (counterAddrTwoStream_valid || counterAddrTwoStream_rValid);
  assign counterAddrTwoStream_s2mPipe_payload = (counterAddrTwoStream_rValid ? counterAddrTwoStream_rData : counterAddrTwoStream_payload);
  always @(*) begin
    counterAddrTwoStream_s2mPipe_ready = counterAddrTwoStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_7) begin
      counterAddrTwoStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_7 = (! counterAddrTwoStream_s2mPipe_m2sPipe_valid);
  assign counterAddrTwoStream_s2mPipe_m2sPipe_valid = counterAddrTwoStream_s2mPipe_rValid;
  assign counterAddrTwoStream_s2mPipe_m2sPipe_payload = counterAddrTwoStream_s2mPipe_rData;
  assign counterAddrTwoStream_s2mPipe_m2sPipe_ready = ((! CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready) || CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready = CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_counterTwoPixelStream_payload = CICC1851_lineBufferTwo_port2;
  assign CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_4 = readStage_counterTwoPixelStream_ready;
    if(when_Stream_l368_8) begin
      CICC1851_4 = 1'b1;
    end
  end

  assign when_Stream_l368_8 = (! readStage_counterTwoPixelStream_valid);
  assign readStage_counterTwoPixelStream_valid = CICC1851_readStage_counterTwoPixelStream_valid;
  assign readStage_counterTwoPixelStream_payload = CICC1851_readStage_counterTwoPixelStream_payload_2;
  assign oddAddrStream_ready = (! oddAddrStream_rValid);
  assign oddAddrStream_s2mPipe_valid = (oddAddrStream_valid || oddAddrStream_rValid);
  assign oddAddrStream_s2mPipe_payload = (oddAddrStream_rValid ? oddAddrStream_rData : oddAddrStream_payload);
  always @(*) begin
    oddAddrStream_s2mPipe_ready = oddAddrStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_9) begin
      oddAddrStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_9 = (! oddAddrStream_s2mPipe_m2sPipe_valid);
  assign oddAddrStream_s2mPipe_m2sPipe_valid = oddAddrStream_s2mPipe_rValid;
  assign oddAddrStream_s2mPipe_m2sPipe_payload = oddAddrStream_s2mPipe_rData;
  assign oddAddrStream_s2mPipe_m2sPipe_ready = ((! CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready) || CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready = CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_oddRowPixelStream_payload = CICC1851_lineBufferOdd_port1;
  assign CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_5 = readStage_oddRowPixelStream_ready;
    if(when_Stream_l368_10) begin
      CICC1851_5 = 1'b1;
    end
  end

  assign when_Stream_l368_10 = (! readStage_oddRowPixelStream_valid);
  assign readStage_oddRowPixelStream_valid = CICC1851_readStage_oddRowPixelStream_valid;
  assign readStage_oddRowPixelStream_payload = CICC1851_readStage_oddRowPixelStream_payload_2;
  assign controlStream_ready = (! controlStream_rValid);
  assign controlStream_s2mPipe_valid = (controlStream_valid || controlStream_rValid);
  assign controlStream_s2mPipe_payload_frameStart = (controlStream_rValid ? controlStream_rData_frameStart : controlStream_payload_frameStart);
  assign controlStream_s2mPipe_payload_rowEnd = (controlStream_rValid ? controlStream_rData_rowEnd : controlStream_payload_rowEnd);
  assign controlStream_s2mPipe_payload_passMode = (controlStream_rValid ? controlStream_rData_passMode : controlStream_payload_passMode);
  assign controlStream_s2mPipe_payload_passValid = (controlStream_rValid ? controlStream_rData_passValid : controlStream_payload_passValid);
  assign controlStream_s2mPipe_payload_onceMode = (controlStream_rValid ? controlStream_rData_onceMode : controlStream_payload_onceMode);
  assign controlStream_s2mPipe_payload_onceValid = (controlStream_rValid ? controlStream_rData_onceValid : controlStream_payload_onceValid);
  assign controlStream_s2mPipe_payload_mainCompare = (controlStream_rValid ? controlStream_rData_mainCompare : controlStream_payload_mainCompare);
  assign controlStream_s2mPipe_payload_counterCompare = (controlStream_rValid ? controlStream_rData_counterCompare : controlStream_payload_counterCompare);
  assign controlStream_s2mPipe_payload_mainDiff = (controlStream_rValid ? controlStream_rData_mainDiff : controlStream_payload_mainDiff);
  assign controlStream_s2mPipe_payload_counterDiff = (controlStream_rValid ? controlStream_rData_counterDiff : controlStream_payload_counterDiff);
  assign controlStream_s2mPipe_payload_twiceCompValid = (controlStream_rValid ? controlStream_rData_twiceCompValid : controlStream_payload_twiceCompValid);
  assign controlStream_s2mPipe_payload_twiceMode = (controlStream_rValid ? controlStream_rData_twiceMode : controlStream_payload_twiceMode);
  assign controlStream_s2mPipe_payload_inpValidFlag = (controlStream_rValid ? controlStream_rData_inpValidFlag : controlStream_payload_inpValidFlag);
  assign controlStream_s2mPipe_payload_oddValid = (controlStream_rValid ? controlStream_rData_oddValid : controlStream_payload_oddValid);
  always @(*) begin
    controlStream_s2mPipe_ready = controlStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_11) begin
      controlStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_11 = (! controlStream_s2mPipe_m2sPipe_valid);
  assign controlStream_s2mPipe_m2sPipe_valid = controlStream_s2mPipe_rValid;
  assign controlStream_s2mPipe_m2sPipe_payload_frameStart = controlStream_s2mPipe_rData_frameStart;
  assign controlStream_s2mPipe_m2sPipe_payload_rowEnd = controlStream_s2mPipe_rData_rowEnd;
  assign controlStream_s2mPipe_m2sPipe_payload_passMode = controlStream_s2mPipe_rData_passMode;
  assign controlStream_s2mPipe_m2sPipe_payload_passValid = controlStream_s2mPipe_rData_passValid;
  assign controlStream_s2mPipe_m2sPipe_payload_onceMode = controlStream_s2mPipe_rData_onceMode;
  assign controlStream_s2mPipe_m2sPipe_payload_onceValid = controlStream_s2mPipe_rData_onceValid;
  assign controlStream_s2mPipe_m2sPipe_payload_mainCompare = controlStream_s2mPipe_rData_mainCompare;
  assign controlStream_s2mPipe_m2sPipe_payload_counterCompare = controlStream_s2mPipe_rData_counterCompare;
  assign controlStream_s2mPipe_m2sPipe_payload_mainDiff = controlStream_s2mPipe_rData_mainDiff;
  assign controlStream_s2mPipe_m2sPipe_payload_counterDiff = controlStream_s2mPipe_rData_counterDiff;
  assign controlStream_s2mPipe_m2sPipe_payload_twiceCompValid = controlStream_s2mPipe_rData_twiceCompValid;
  assign controlStream_s2mPipe_m2sPipe_payload_twiceMode = controlStream_s2mPipe_rData_twiceMode;
  assign controlStream_s2mPipe_m2sPipe_payload_inpValidFlag = controlStream_s2mPipe_rData_inpValidFlag;
  assign controlStream_s2mPipe_m2sPipe_payload_oddValid = controlStream_s2mPipe_rData_oddValid;
  always @(*) begin
    controlStream_s2mPipe_m2sPipe_ready = controlStream_s2mPipe_m2sPipe_m2sPipe_ready;
    if(when_Stream_l368_12) begin
      controlStream_s2mPipe_m2sPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_12 = (! controlStream_s2mPipe_m2sPipe_m2sPipe_valid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_valid = controlStream_s2mPipe_m2sPipe_rValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_frameStart = controlStream_s2mPipe_m2sPipe_rData_frameStart;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_rowEnd = controlStream_s2mPipe_m2sPipe_rData_rowEnd;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passMode = controlStream_s2mPipe_m2sPipe_rData_passMode;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passValid = controlStream_s2mPipe_m2sPipe_rData_passValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceMode = controlStream_s2mPipe_m2sPipe_rData_onceMode;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceValid = controlStream_s2mPipe_m2sPipe_rData_onceValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainCompare = controlStream_s2mPipe_m2sPipe_rData_mainCompare;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterCompare = controlStream_s2mPipe_m2sPipe_rData_counterCompare;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDiff = controlStream_s2mPipe_m2sPipe_rData_mainDiff;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDiff = controlStream_s2mPipe_m2sPipe_rData_counterDiff;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceCompValid = controlStream_s2mPipe_m2sPipe_rData_twiceCompValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceMode = controlStream_s2mPipe_m2sPipe_rData_twiceMode;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_inpValidFlag = controlStream_s2mPipe_m2sPipe_rData_inpValidFlag;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_oddValid = controlStream_s2mPipe_m2sPipe_rData_oddValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_ready = (! controlStream_s2mPipe_m2sPipe_m2sPipe_rValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_valid = (controlStream_s2mPipe_m2sPipe_m2sPipe_valid || controlStream_s2mPipe_m2sPipe_m2sPipe_rValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_frameStart = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_frameStart : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_frameStart);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_rowEnd = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_rowEnd : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_rowEnd);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_passMode = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_passMode : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passMode);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_passValid = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_passValid : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_onceMode = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_onceMode : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceMode);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_onceValid = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_onceValid : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainCompare = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainCompare : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainCompare);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterCompare = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterCompare : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterCompare);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainDiff = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainDiff : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDiff);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterDiff = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterDiff : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDiff);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_twiceCompValid = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_twiceCompValid : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceCompValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_twiceMode = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_twiceMode : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceMode);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_inpValidFlag = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_inpValidFlag : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_inpValidFlag);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_oddValid = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_oddValid : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_oddValid);
  always @(*) begin
    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready = readStage_controlPipe_ready;
    if(when_Stream_l368_13) begin
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_13 = (! readStage_controlPipe_valid);
  assign readStage_controlPipe_valid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rValid;
  assign readStage_controlPipe_payload_frameStart = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_frameStart;
  assign readStage_controlPipe_payload_rowEnd = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_rowEnd;
  assign readStage_controlPipe_payload_passMode = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_passMode;
  assign readStage_controlPipe_payload_passValid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_passValid;
  assign readStage_controlPipe_payload_onceMode = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_onceMode;
  assign readStage_controlPipe_payload_onceValid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_onceValid;
  assign readStage_controlPipe_payload_mainCompare = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainCompare;
  assign readStage_controlPipe_payload_counterCompare = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterCompare;
  assign readStage_controlPipe_payload_mainDiff = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainDiff;
  assign readStage_controlPipe_payload_counterDiff = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterDiff;
  assign readStage_controlPipe_payload_twiceCompValid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_twiceCompValid;
  assign readStage_controlPipe_payload_twiceMode = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_twiceMode;
  assign readStage_controlPipe_payload_inpValidFlag = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_inpValidFlag;
  assign readStage_controlPipe_payload_oddValid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_oddValid;
  assign readStage_mainOnePixelStream_ready = (! readStage_mainOnePixelStream_rValid);
  assign readStage_mainOnePixelStream_s2mPipe_valid = (readStage_mainOnePixelStream_valid || readStage_mainOnePixelStream_rValid);
  assign readStage_mainOnePixelStream_s2mPipe_payload = (readStage_mainOnePixelStream_rValid ? readStage_mainOnePixelStream_rData : readStage_mainOnePixelStream_payload);
  always @(*) begin
    readStage_mainOnePixelStream_s2mPipe_ready = compareStage_mainOnePixelStream_ready;
    if(when_Stream_l368_14) begin
      readStage_mainOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_14 = (! compareStage_mainOnePixelStream_valid);
  assign compareStage_mainOnePixelStream_valid = readStage_mainOnePixelStream_s2mPipe_rValid;
  assign compareStage_mainOnePixelStream_payload = readStage_mainOnePixelStream_s2mPipe_rData;
  assign readStage_counterOnePixelStream_ready = (! readStage_counterOnePixelStream_rValid);
  assign readStage_counterOnePixelStream_s2mPipe_valid = (readStage_counterOnePixelStream_valid || readStage_counterOnePixelStream_rValid);
  assign readStage_counterOnePixelStream_s2mPipe_payload = (readStage_counterOnePixelStream_rValid ? readStage_counterOnePixelStream_rData : readStage_counterOnePixelStream_payload);
  always @(*) begin
    readStage_counterOnePixelStream_s2mPipe_ready = compareStage_counterOnePixelStream_ready;
    if(when_Stream_l368_15) begin
      readStage_counterOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_15 = (! compareStage_counterOnePixelStream_valid);
  assign compareStage_counterOnePixelStream_valid = readStage_counterOnePixelStream_s2mPipe_rValid;
  assign compareStage_counterOnePixelStream_payload = readStage_counterOnePixelStream_s2mPipe_rData;
  assign readStage_mainTwoPixelStream_ready = (! readStage_mainTwoPixelStream_rValid);
  assign readStage_mainTwoPixelStream_s2mPipe_valid = (readStage_mainTwoPixelStream_valid || readStage_mainTwoPixelStream_rValid);
  assign readStage_mainTwoPixelStream_s2mPipe_payload = (readStage_mainTwoPixelStream_rValid ? readStage_mainTwoPixelStream_rData : readStage_mainTwoPixelStream_payload);
  always @(*) begin
    readStage_mainTwoPixelStream_s2mPipe_ready = compareStage_mainTwoPixelStream_ready;
    if(when_Stream_l368_16) begin
      readStage_mainTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_16 = (! compareStage_mainTwoPixelStream_valid);
  assign compareStage_mainTwoPixelStream_valid = readStage_mainTwoPixelStream_s2mPipe_rValid;
  assign compareStage_mainTwoPixelStream_payload = readStage_mainTwoPixelStream_s2mPipe_rData;
  assign readStage_counterTwoPixelStream_ready = (! readStage_counterTwoPixelStream_rValid);
  assign readStage_counterTwoPixelStream_s2mPipe_valid = (readStage_counterTwoPixelStream_valid || readStage_counterTwoPixelStream_rValid);
  assign readStage_counterTwoPixelStream_s2mPipe_payload = (readStage_counterTwoPixelStream_rValid ? readStage_counterTwoPixelStream_rData : readStage_counterTwoPixelStream_payload);
  always @(*) begin
    readStage_counterTwoPixelStream_s2mPipe_ready = compareStage_counterTwoPixelStream_ready;
    if(when_Stream_l368_17) begin
      readStage_counterTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_17 = (! compareStage_counterTwoPixelStream_valid);
  assign compareStage_counterTwoPixelStream_valid = readStage_counterTwoPixelStream_s2mPipe_rValid;
  assign compareStage_counterTwoPixelStream_payload = readStage_counterTwoPixelStream_s2mPipe_rData;
  assign readStage_oddRowPixelStream_ready = (! readStage_oddRowPixelStream_rValid);
  assign readStage_oddRowPixelStream_s2mPipe_valid = (readStage_oddRowPixelStream_valid || readStage_oddRowPixelStream_rValid);
  assign readStage_oddRowPixelStream_s2mPipe_payload = (readStage_oddRowPixelStream_rValid ? readStage_oddRowPixelStream_rData : readStage_oddRowPixelStream_payload);
  always @(*) begin
    readStage_oddRowPixelStream_s2mPipe_ready = compareStage_oddRowPixelStream_ready;
    if(when_Stream_l368_18) begin
      readStage_oddRowPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_18 = (! compareStage_oddRowPixelStream_valid);
  assign compareStage_oddRowPixelStream_valid = readStage_oddRowPixelStream_s2mPipe_rValid;
  assign compareStage_oddRowPixelStream_payload = readStage_oddRowPixelStream_s2mPipe_rData;
  always @(*) begin
    CICC1851_readStage_controlPipe_translated_payload_mainCompare = readStage_controlPipe_payload_mainCompare;
    if(readStage_controlPipe_payload_onceValid) begin
      case(readStage_controlPipe_payload_onceMode)
        3'b000 : begin
          if(when_SuperResolutionPart2_l290) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        3'b001 : begin
          if(when_SuperResolutionPart2_l294) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        3'b010 : begin
          if(when_SuperResolutionPart2_l298) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        3'b011 : begin
          if(when_SuperResolutionPart2_l302) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        3'b100 : begin
          CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
        end
        3'b101 : begin
          CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
        end
        default : begin
        end
      endcase
    end
    if(readStage_controlPipe_payload_twiceCompValid) begin
      case(readStage_controlPipe_payload_twiceMode)
        3'b000 : begin
          if(when_SuperResolutionPart2_l313) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        3'b001 : begin
          if(when_SuperResolutionPart2_l319) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        3'b010 : begin
          CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
        end
        3'b011 : begin
          if(when_SuperResolutionPart2_l326) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        3'b100 : begin
          CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
        end
        3'b101 : begin
          if(when_SuperResolutionPart2_l331) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    CICC1851_readStage_controlPipe_translated_payload_counterCompare = readStage_controlPipe_payload_counterCompare;
    if(readStage_controlPipe_payload_twiceCompValid) begin
      case(readStage_controlPipe_payload_twiceMode)
        3'b000 : begin
          if(when_SuperResolutionPart2_l315) begin
            CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
          end
        end
        3'b001 : begin
          if(when_SuperResolutionPart2_l321) begin
            CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
          end
        end
        default : begin
        end
      endcase
    end
  end

  assign when_SuperResolutionPart2_l290 = (readStage_counterOnePixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart2_l294 = (readStage_counterTwoPixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart2_l298 = (readStage_mainTwoPixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart2_l302 = (readStage_mainOnePixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart2_l313 = (readStage_mainTwoPixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart2_l315 = (readStage_counterOnePixelStream_payload <= readStage_counterTwoPixelStream_payload);
  assign when_SuperResolutionPart2_l319 = (readStage_mainOnePixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart2_l321 = (readStage_counterTwoPixelStream_payload <= readStage_counterOnePixelStream_payload);
  assign when_SuperResolutionPart2_l326 = (readStage_counterTwoPixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart2_l331 = (readStage_counterOnePixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign readStage_controlPipe_translated_valid = readStage_controlPipe_valid;
  assign readStage_controlPipe_ready = readStage_controlPipe_translated_ready;
  assign readStage_controlPipe_translated_payload_frameStart = readStage_controlPipe_payload_frameStart;
  assign readStage_controlPipe_translated_payload_rowEnd = readStage_controlPipe_payload_rowEnd;
  assign readStage_controlPipe_translated_payload_passMode = readStage_controlPipe_payload_passMode;
  assign readStage_controlPipe_translated_payload_passValid = readStage_controlPipe_payload_passValid;
  assign readStage_controlPipe_translated_payload_onceMode = readStage_controlPipe_payload_onceMode;
  assign readStage_controlPipe_translated_payload_onceValid = readStage_controlPipe_payload_onceValid;
  assign readStage_controlPipe_translated_payload_mainCompare = CICC1851_readStage_controlPipe_translated_payload_mainCompare;
  assign readStage_controlPipe_translated_payload_counterCompare = CICC1851_readStage_controlPipe_translated_payload_counterCompare;
  assign readStage_controlPipe_translated_payload_mainDiff = readStage_controlPipe_payload_mainDiff;
  assign readStage_controlPipe_translated_payload_counterDiff = readStage_controlPipe_payload_counterDiff;
  assign readStage_controlPipe_translated_payload_twiceCompValid = readStage_controlPipe_payload_twiceCompValid;
  assign readStage_controlPipe_translated_payload_twiceMode = readStage_controlPipe_payload_twiceMode;
  assign readStage_controlPipe_translated_payload_inpValidFlag = readStage_controlPipe_payload_inpValidFlag;
  assign readStage_controlPipe_translated_payload_oddValid = readStage_controlPipe_payload_oddValid;
  assign readStage_controlPipe_translated_ready = (! readStage_controlPipe_translated_rValid);
  assign readStage_controlPipe_translated_s2mPipe_valid = (readStage_controlPipe_translated_valid || readStage_controlPipe_translated_rValid);
  assign readStage_controlPipe_translated_s2mPipe_payload_frameStart = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_frameStart : readStage_controlPipe_translated_payload_frameStart);
  assign readStage_controlPipe_translated_s2mPipe_payload_rowEnd = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_rowEnd : readStage_controlPipe_translated_payload_rowEnd);
  assign readStage_controlPipe_translated_s2mPipe_payload_passMode = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_passMode : readStage_controlPipe_translated_payload_passMode);
  assign readStage_controlPipe_translated_s2mPipe_payload_passValid = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_passValid : readStage_controlPipe_translated_payload_passValid);
  assign readStage_controlPipe_translated_s2mPipe_payload_onceMode = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_onceMode : readStage_controlPipe_translated_payload_onceMode);
  assign readStage_controlPipe_translated_s2mPipe_payload_onceValid = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_onceValid : readStage_controlPipe_translated_payload_onceValid);
  assign readStage_controlPipe_translated_s2mPipe_payload_mainCompare = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_mainCompare : readStage_controlPipe_translated_payload_mainCompare);
  assign readStage_controlPipe_translated_s2mPipe_payload_counterCompare = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_counterCompare : readStage_controlPipe_translated_payload_counterCompare);
  assign readStage_controlPipe_translated_s2mPipe_payload_mainDiff = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_mainDiff : readStage_controlPipe_translated_payload_mainDiff);
  assign readStage_controlPipe_translated_s2mPipe_payload_counterDiff = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_counterDiff : readStage_controlPipe_translated_payload_counterDiff);
  assign readStage_controlPipe_translated_s2mPipe_payload_twiceCompValid = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_twiceCompValid : readStage_controlPipe_translated_payload_twiceCompValid);
  assign readStage_controlPipe_translated_s2mPipe_payload_twiceMode = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_twiceMode : readStage_controlPipe_translated_payload_twiceMode);
  assign readStage_controlPipe_translated_s2mPipe_payload_inpValidFlag = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_inpValidFlag : readStage_controlPipe_translated_payload_inpValidFlag);
  assign readStage_controlPipe_translated_s2mPipe_payload_oddValid = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_oddValid : readStage_controlPipe_translated_payload_oddValid);
  always @(*) begin
    readStage_controlPipe_translated_s2mPipe_ready = compareStage_controlPipe_ready;
    if(when_Stream_l368_19) begin
      readStage_controlPipe_translated_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_19 = (! compareStage_controlPipe_valid);
  assign compareStage_controlPipe_valid = readStage_controlPipe_translated_s2mPipe_rValid;
  assign compareStage_controlPipe_payload_frameStart = readStage_controlPipe_translated_s2mPipe_rData_frameStart;
  assign compareStage_controlPipe_payload_rowEnd = readStage_controlPipe_translated_s2mPipe_rData_rowEnd;
  assign compareStage_controlPipe_payload_passMode = readStage_controlPipe_translated_s2mPipe_rData_passMode;
  assign compareStage_controlPipe_payload_passValid = readStage_controlPipe_translated_s2mPipe_rData_passValid;
  assign compareStage_controlPipe_payload_onceMode = readStage_controlPipe_translated_s2mPipe_rData_onceMode;
  assign compareStage_controlPipe_payload_onceValid = readStage_controlPipe_translated_s2mPipe_rData_onceValid;
  assign compareStage_controlPipe_payload_mainCompare = readStage_controlPipe_translated_s2mPipe_rData_mainCompare;
  assign compareStage_controlPipe_payload_counterCompare = readStage_controlPipe_translated_s2mPipe_rData_counterCompare;
  assign compareStage_controlPipe_payload_mainDiff = readStage_controlPipe_translated_s2mPipe_rData_mainDiff;
  assign compareStage_controlPipe_payload_counterDiff = readStage_controlPipe_translated_s2mPipe_rData_counterDiff;
  assign compareStage_controlPipe_payload_twiceCompValid = readStage_controlPipe_translated_s2mPipe_rData_twiceCompValid;
  assign compareStage_controlPipe_payload_twiceMode = readStage_controlPipe_translated_s2mPipe_rData_twiceMode;
  assign compareStage_controlPipe_payload_inpValidFlag = readStage_controlPipe_translated_s2mPipe_rData_inpValidFlag;
  assign compareStage_controlPipe_payload_oddValid = readStage_controlPipe_translated_s2mPipe_rData_oddValid;
  assign compareStage_mainOnePixelStream_ready = (! compareStage_mainOnePixelStream_rValid);
  assign compareStage_mainOnePixelStream_s2mPipe_valid = (compareStage_mainOnePixelStream_valid || compareStage_mainOnePixelStream_rValid);
  assign compareStage_mainOnePixelStream_s2mPipe_payload = (compareStage_mainOnePixelStream_rValid ? compareStage_mainOnePixelStream_rData : compareStage_mainOnePixelStream_payload);
  always @(*) begin
    compareStage_mainOnePixelStream_s2mPipe_ready = diffStage_mainOnePixelStream_ready;
    if(when_Stream_l368_20) begin
      compareStage_mainOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_20 = (! diffStage_mainOnePixelStream_valid);
  assign diffStage_mainOnePixelStream_valid = compareStage_mainOnePixelStream_s2mPipe_rValid;
  assign diffStage_mainOnePixelStream_payload = compareStage_mainOnePixelStream_s2mPipe_rData;
  assign compareStage_counterOnePixelStream_ready = (! compareStage_counterOnePixelStream_rValid);
  assign compareStage_counterOnePixelStream_s2mPipe_valid = (compareStage_counterOnePixelStream_valid || compareStage_counterOnePixelStream_rValid);
  assign compareStage_counterOnePixelStream_s2mPipe_payload = (compareStage_counterOnePixelStream_rValid ? compareStage_counterOnePixelStream_rData : compareStage_counterOnePixelStream_payload);
  always @(*) begin
    compareStage_counterOnePixelStream_s2mPipe_ready = diffStage_counterOnePixelStream_ready;
    if(when_Stream_l368_21) begin
      compareStage_counterOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_21 = (! diffStage_counterOnePixelStream_valid);
  assign diffStage_counterOnePixelStream_valid = compareStage_counterOnePixelStream_s2mPipe_rValid;
  assign diffStage_counterOnePixelStream_payload = compareStage_counterOnePixelStream_s2mPipe_rData;
  assign compareStage_mainTwoPixelStream_ready = (! compareStage_mainTwoPixelStream_rValid);
  assign compareStage_mainTwoPixelStream_s2mPipe_valid = (compareStage_mainTwoPixelStream_valid || compareStage_mainTwoPixelStream_rValid);
  assign compareStage_mainTwoPixelStream_s2mPipe_payload = (compareStage_mainTwoPixelStream_rValid ? compareStage_mainTwoPixelStream_rData : compareStage_mainTwoPixelStream_payload);
  always @(*) begin
    compareStage_mainTwoPixelStream_s2mPipe_ready = diffStage_mainTwoPixelStream_ready;
    if(when_Stream_l368_22) begin
      compareStage_mainTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_22 = (! diffStage_mainTwoPixelStream_valid);
  assign diffStage_mainTwoPixelStream_valid = compareStage_mainTwoPixelStream_s2mPipe_rValid;
  assign diffStage_mainTwoPixelStream_payload = compareStage_mainTwoPixelStream_s2mPipe_rData;
  assign compareStage_counterTwoPixelStream_ready = (! compareStage_counterTwoPixelStream_rValid);
  assign compareStage_counterTwoPixelStream_s2mPipe_valid = (compareStage_counterTwoPixelStream_valid || compareStage_counterTwoPixelStream_rValid);
  assign compareStage_counterTwoPixelStream_s2mPipe_payload = (compareStage_counterTwoPixelStream_rValid ? compareStage_counterTwoPixelStream_rData : compareStage_counterTwoPixelStream_payload);
  always @(*) begin
    compareStage_counterTwoPixelStream_s2mPipe_ready = diffStage_counterTwoPixelStream_ready;
    if(when_Stream_l368_23) begin
      compareStage_counterTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_23 = (! diffStage_counterTwoPixelStream_valid);
  assign diffStage_counterTwoPixelStream_valid = compareStage_counterTwoPixelStream_s2mPipe_rValid;
  assign diffStage_counterTwoPixelStream_payload = compareStage_counterTwoPixelStream_s2mPipe_rData;
  assign compareStage_oddRowPixelStream_ready = (! compareStage_oddRowPixelStream_rValid);
  assign compareStage_oddRowPixelStream_s2mPipe_valid = (compareStage_oddRowPixelStream_valid || compareStage_oddRowPixelStream_rValid);
  assign compareStage_oddRowPixelStream_s2mPipe_payload = (compareStage_oddRowPixelStream_rValid ? compareStage_oddRowPixelStream_rData : compareStage_oddRowPixelStream_payload);
  always @(*) begin
    compareStage_oddRowPixelStream_s2mPipe_ready = diffStage_oddRowPixelStream_ready;
    if(when_Stream_l368_24) begin
      compareStage_oddRowPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_24 = (! diffStage_oddRowPixelStream_valid);
  assign diffStage_oddRowPixelStream_valid = compareStage_oddRowPixelStream_s2mPipe_rValid;
  assign diffStage_oddRowPixelStream_payload = compareStage_oddRowPixelStream_s2mPipe_rData;
  always @(*) begin
    CICC1851_compareStage_controlPipe_translated_payload_mainDiff = compareStage_controlPipe_payload_mainDiff;
    if(compareStage_controlPipe_payload_onceValid) begin
      case(compareStage_controlPipe_payload_onceMode)
        3'b000 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_counterOnePixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterOnePixelStream_payload - compareStage_mainOnePixelStream_payload);
          end
        end
        3'b001 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterTwoPixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainTwoPixelStream_payload);
          end
        end
        3'b010 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_mainTwoPixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_mainOnePixelStream_payload);
          end
        end
        3'b011 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_mainOnePixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_mainTwoPixelStream_payload);
          end
        end
        3'b100 : begin
          CICC1851_compareStage_controlPipe_translated_payload_mainDiff = 8'h0;
        end
        3'b101 : begin
          CICC1851_compareStage_controlPipe_translated_payload_mainDiff = 8'h0;
        end
        default : begin
        end
      endcase
    end
    if(compareStage_controlPipe_payload_twiceCompValid) begin
      case(compareStage_controlPipe_payload_twiceMode)
        3'b000 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_mainTwoPixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_mainOnePixelStream_payload);
          end
        end
        3'b001 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_mainOnePixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_mainTwoPixelStream_payload);
          end
        end
        3'b010 : begin
          CICC1851_compareStage_controlPipe_translated_payload_mainDiff = 8'h0;
        end
        3'b011 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterTwoPixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainTwoPixelStream_payload);
          end
        end
        3'b100 : begin
          CICC1851_compareStage_controlPipe_translated_payload_mainDiff = 8'h0;
        end
        3'b101 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_counterOnePixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterOnePixelStream_payload - compareStage_mainOnePixelStream_payload);
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    CICC1851_compareStage_controlPipe_translated_payload_counterDiff = compareStage_controlPipe_payload_counterDiff;
    if(compareStage_controlPipe_payload_twiceCompValid) begin
      case(compareStage_controlPipe_payload_twiceMode)
        3'b000 : begin
          if(compareStage_controlPipe_payload_counterCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterTwoPixelStream_payload - compareStage_counterOnePixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterOnePixelStream_payload - compareStage_counterTwoPixelStream_payload);
          end
        end
        3'b001 : begin
          if(compareStage_controlPipe_payload_counterCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterOnePixelStream_payload - compareStage_counterTwoPixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterTwoPixelStream_payload - compareStage_counterOnePixelStream_payload);
          end
        end
        default : begin
        end
      endcase
    end
  end

  assign compareStage_controlPipe_translated_valid = compareStage_controlPipe_valid;
  assign compareStage_controlPipe_ready = compareStage_controlPipe_translated_ready;
  assign compareStage_controlPipe_translated_payload_frameStart = compareStage_controlPipe_payload_frameStart;
  assign compareStage_controlPipe_translated_payload_rowEnd = compareStage_controlPipe_payload_rowEnd;
  assign compareStage_controlPipe_translated_payload_passMode = compareStage_controlPipe_payload_passMode;
  assign compareStage_controlPipe_translated_payload_passValid = compareStage_controlPipe_payload_passValid;
  assign compareStage_controlPipe_translated_payload_onceMode = compareStage_controlPipe_payload_onceMode;
  assign compareStage_controlPipe_translated_payload_onceValid = compareStage_controlPipe_payload_onceValid;
  assign compareStage_controlPipe_translated_payload_mainCompare = compareStage_controlPipe_payload_mainCompare;
  assign compareStage_controlPipe_translated_payload_counterCompare = compareStage_controlPipe_payload_counterCompare;
  assign compareStage_controlPipe_translated_payload_mainDiff = CICC1851_compareStage_controlPipe_translated_payload_mainDiff;
  assign compareStage_controlPipe_translated_payload_counterDiff = CICC1851_compareStage_controlPipe_translated_payload_counterDiff;
  assign compareStage_controlPipe_translated_payload_twiceCompValid = compareStage_controlPipe_payload_twiceCompValid;
  assign compareStage_controlPipe_translated_payload_twiceMode = compareStage_controlPipe_payload_twiceMode;
  assign compareStage_controlPipe_translated_payload_inpValidFlag = compareStage_controlPipe_payload_inpValidFlag;
  assign compareStage_controlPipe_translated_payload_oddValid = compareStage_controlPipe_payload_oddValid;
  assign compareStage_controlPipe_translated_ready = (! compareStage_controlPipe_translated_rValid);
  assign compareStage_controlPipe_translated_s2mPipe_valid = (compareStage_controlPipe_translated_valid || compareStage_controlPipe_translated_rValid);
  assign compareStage_controlPipe_translated_s2mPipe_payload_frameStart = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_frameStart : compareStage_controlPipe_translated_payload_frameStart);
  assign compareStage_controlPipe_translated_s2mPipe_payload_rowEnd = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_rowEnd : compareStage_controlPipe_translated_payload_rowEnd);
  assign compareStage_controlPipe_translated_s2mPipe_payload_passMode = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_passMode : compareStage_controlPipe_translated_payload_passMode);
  assign compareStage_controlPipe_translated_s2mPipe_payload_passValid = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_passValid : compareStage_controlPipe_translated_payload_passValid);
  assign compareStage_controlPipe_translated_s2mPipe_payload_onceMode = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_onceMode : compareStage_controlPipe_translated_payload_onceMode);
  assign compareStage_controlPipe_translated_s2mPipe_payload_onceValid = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_onceValid : compareStage_controlPipe_translated_payload_onceValid);
  assign compareStage_controlPipe_translated_s2mPipe_payload_mainCompare = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_mainCompare : compareStage_controlPipe_translated_payload_mainCompare);
  assign compareStage_controlPipe_translated_s2mPipe_payload_counterCompare = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_counterCompare : compareStage_controlPipe_translated_payload_counterCompare);
  assign compareStage_controlPipe_translated_s2mPipe_payload_mainDiff = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_mainDiff : compareStage_controlPipe_translated_payload_mainDiff);
  assign compareStage_controlPipe_translated_s2mPipe_payload_counterDiff = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_counterDiff : compareStage_controlPipe_translated_payload_counterDiff);
  assign compareStage_controlPipe_translated_s2mPipe_payload_twiceCompValid = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_twiceCompValid : compareStage_controlPipe_translated_payload_twiceCompValid);
  assign compareStage_controlPipe_translated_s2mPipe_payload_twiceMode = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_twiceMode : compareStage_controlPipe_translated_payload_twiceMode);
  assign compareStage_controlPipe_translated_s2mPipe_payload_inpValidFlag = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_inpValidFlag : compareStage_controlPipe_translated_payload_inpValidFlag);
  assign compareStage_controlPipe_translated_s2mPipe_payload_oddValid = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_oddValid : compareStage_controlPipe_translated_payload_oddValid);
  always @(*) begin
    compareStage_controlPipe_translated_s2mPipe_ready = diffStage_controlPipe_ready;
    if(when_Stream_l368_25) begin
      compareStage_controlPipe_translated_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_25 = (! diffStage_controlPipe_valid);
  assign diffStage_controlPipe_valid = compareStage_controlPipe_translated_s2mPipe_rValid;
  assign diffStage_controlPipe_payload_frameStart = compareStage_controlPipe_translated_s2mPipe_rData_frameStart;
  assign diffStage_controlPipe_payload_rowEnd = compareStage_controlPipe_translated_s2mPipe_rData_rowEnd;
  assign diffStage_controlPipe_payload_passMode = compareStage_controlPipe_translated_s2mPipe_rData_passMode;
  assign diffStage_controlPipe_payload_passValid = compareStage_controlPipe_translated_s2mPipe_rData_passValid;
  assign diffStage_controlPipe_payload_onceMode = compareStage_controlPipe_translated_s2mPipe_rData_onceMode;
  assign diffStage_controlPipe_payload_onceValid = compareStage_controlPipe_translated_s2mPipe_rData_onceValid;
  assign diffStage_controlPipe_payload_mainCompare = compareStage_controlPipe_translated_s2mPipe_rData_mainCompare;
  assign diffStage_controlPipe_payload_counterCompare = compareStage_controlPipe_translated_s2mPipe_rData_counterCompare;
  assign diffStage_controlPipe_payload_mainDiff = compareStage_controlPipe_translated_s2mPipe_rData_mainDiff;
  assign diffStage_controlPipe_payload_counterDiff = compareStage_controlPipe_translated_s2mPipe_rData_counterDiff;
  assign diffStage_controlPipe_payload_twiceCompValid = compareStage_controlPipe_translated_s2mPipe_rData_twiceCompValid;
  assign diffStage_controlPipe_payload_twiceMode = compareStage_controlPipe_translated_s2mPipe_rData_twiceMode;
  assign diffStage_controlPipe_payload_inpValidFlag = compareStage_controlPipe_translated_s2mPipe_rData_inpValidFlag;
  assign diffStage_controlPipe_payload_oddValid = compareStage_controlPipe_translated_s2mPipe_rData_oddValid;
  assign diffStage_mainOnePixelStream_ready = (! diffStage_mainOnePixelStream_rValid);
  assign diffStage_mainOnePixelStream_s2mPipe_valid = (diffStage_mainOnePixelStream_valid || diffStage_mainOnePixelStream_rValid);
  assign diffStage_mainOnePixelStream_s2mPipe_payload = (diffStage_mainOnePixelStream_rValid ? diffStage_mainOnePixelStream_rData : diffStage_mainOnePixelStream_payload);
  always @(*) begin
    diffStage_mainOnePixelStream_s2mPipe_ready = resultStage_mainOnePixelStream_ready;
    if(when_Stream_l368_26) begin
      diffStage_mainOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_26 = (! resultStage_mainOnePixelStream_valid);
  assign resultStage_mainOnePixelStream_valid = diffStage_mainOnePixelStream_s2mPipe_rValid;
  assign resultStage_mainOnePixelStream_payload = diffStage_mainOnePixelStream_s2mPipe_rData;
  assign diffStage_counterOnePixelStream_ready = (! diffStage_counterOnePixelStream_rValid);
  assign diffStage_counterOnePixelStream_s2mPipe_valid = (diffStage_counterOnePixelStream_valid || diffStage_counterOnePixelStream_rValid);
  assign diffStage_counterOnePixelStream_s2mPipe_payload = (diffStage_counterOnePixelStream_rValid ? diffStage_counterOnePixelStream_rData : diffStage_counterOnePixelStream_payload);
  always @(*) begin
    diffStage_counterOnePixelStream_s2mPipe_ready = resultStage_counterOnePixelStream_ready;
    if(when_Stream_l368_27) begin
      diffStage_counterOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_27 = (! resultStage_counterOnePixelStream_valid);
  assign resultStage_counterOnePixelStream_valid = diffStage_counterOnePixelStream_s2mPipe_rValid;
  assign resultStage_counterOnePixelStream_payload = diffStage_counterOnePixelStream_s2mPipe_rData;
  assign diffStage_mainTwoPixelStream_ready = (! diffStage_mainTwoPixelStream_rValid);
  assign diffStage_mainTwoPixelStream_s2mPipe_valid = (diffStage_mainTwoPixelStream_valid || diffStage_mainTwoPixelStream_rValid);
  assign diffStage_mainTwoPixelStream_s2mPipe_payload = (diffStage_mainTwoPixelStream_rValid ? diffStage_mainTwoPixelStream_rData : diffStage_mainTwoPixelStream_payload);
  always @(*) begin
    diffStage_mainTwoPixelStream_s2mPipe_ready = resultStage_mainTwoPixelStream_ready;
    if(when_Stream_l368_28) begin
      diffStage_mainTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_28 = (! resultStage_mainTwoPixelStream_valid);
  assign resultStage_mainTwoPixelStream_valid = diffStage_mainTwoPixelStream_s2mPipe_rValid;
  assign resultStage_mainTwoPixelStream_payload = diffStage_mainTwoPixelStream_s2mPipe_rData;
  assign diffStage_counterTwoPixelStream_ready = (! diffStage_counterTwoPixelStream_rValid);
  assign diffStage_counterTwoPixelStream_s2mPipe_valid = (diffStage_counterTwoPixelStream_valid || diffStage_counterTwoPixelStream_rValid);
  assign diffStage_counterTwoPixelStream_s2mPipe_payload = (diffStage_counterTwoPixelStream_rValid ? diffStage_counterTwoPixelStream_rData : diffStage_counterTwoPixelStream_payload);
  always @(*) begin
    diffStage_counterTwoPixelStream_s2mPipe_ready = resultStage_counterTwoPixelStream_ready;
    if(when_Stream_l368_29) begin
      diffStage_counterTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_29 = (! resultStage_counterTwoPixelStream_valid);
  assign resultStage_counterTwoPixelStream_valid = diffStage_counterTwoPixelStream_s2mPipe_rValid;
  assign resultStage_counterTwoPixelStream_payload = diffStage_counterTwoPixelStream_s2mPipe_rData;
  assign diffStage_oddRowPixelStream_ready = (! diffStage_oddRowPixelStream_rValid);
  assign diffStage_oddRowPixelStream_s2mPipe_valid = (diffStage_oddRowPixelStream_valid || diffStage_oddRowPixelStream_rValid);
  assign diffStage_oddRowPixelStream_s2mPipe_payload = (diffStage_oddRowPixelStream_rValid ? diffStage_oddRowPixelStream_rData : diffStage_oddRowPixelStream_payload);
  always @(*) begin
    diffStage_oddRowPixelStream_s2mPipe_ready = resultStage_oddRowPixelStream_ready;
    if(when_Stream_l368_30) begin
      diffStage_oddRowPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_30 = (! resultStage_oddRowPixelStream_valid);
  assign resultStage_oddRowPixelStream_valid = diffStage_oddRowPixelStream_s2mPipe_rValid;
  assign resultStage_oddRowPixelStream_payload = diffStage_oddRowPixelStream_s2mPipe_rData;
  assign diffStage_controlPipe_ready = diffStage_controlPipe_fork_io_input_ready;
  assign CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceMode = diffStage_controlPipe_payload_onceMode;
  assign CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceValid = diffStage_controlPipe_payload_onceValid;
  assign CICC1851_when_SuperResolutionPart2_l419 = diffStage_controlPipe_payload_mainDiff;
  assign CICC1851_when_SuperResolutionPart2_l428 = diffStage_controlPipe_payload_counterDiff;
  assign CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceCompValid = diffStage_controlPipe_payload_twiceCompValid;
  assign CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceMode = diffStage_controlPipe_payload_twiceMode;
  always @(*) begin
    CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag = diffStage_controlPipe_payload_inpValidFlag;
    if(CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceValid) begin
      case(CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceMode)
        3'b000 : begin
          if(when_SuperResolutionPart2_l419) begin
            CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag = 1'b0;
          end
        end
        3'b001 : begin
          if(when_SuperResolutionPart2_l420) begin
            CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag = 1'b0;
          end
        end
        3'b010 : begin
          if(when_SuperResolutionPart2_l421) begin
            CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag = 1'b0;
          end
        end
        3'b011 : begin
          if(when_SuperResolutionPart2_l422) begin
            CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag = 1'b0;
          end
        end
        default : begin
        end
      endcase
    end
    if(CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceCompValid) begin
      case(CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceMode)
        3'b000 : begin
          if(when_SuperResolutionPart2_l428) begin
            CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag = 1'b0;
          end
        end
        3'b001 : begin
          if(when_SuperResolutionPart2_l429) begin
            CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag = 1'b0;
          end
        end
        3'b011 : begin
          if(when_SuperResolutionPart2_l430) begin
            CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag = 1'b0;
          end
        end
        3'b101 : begin
          if(when_SuperResolutionPart2_l431) begin
            CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag = 1'b0;
          end
        end
        default : begin
        end
      endcase
    end
  end

  assign when_SuperResolutionPart2_l419 = (inpThreshold <= CICC1851_when_SuperResolutionPart2_l419);
  assign when_SuperResolutionPart2_l420 = (inpThreshold <= CICC1851_when_SuperResolutionPart2_l419);
  assign when_SuperResolutionPart2_l421 = (inpThreshold <= CICC1851_when_SuperResolutionPart2_l419);
  assign when_SuperResolutionPart2_l422 = (inpThreshold <= CICC1851_when_SuperResolutionPart2_l419);
  assign when_SuperResolutionPart2_l428 = ((inpThreshold <= CICC1851_when_SuperResolutionPart2_l419) && (inpThreshold <= CICC1851_when_SuperResolutionPart2_l428));
  assign when_SuperResolutionPart2_l429 = ((inpThreshold <= CICC1851_when_SuperResolutionPart2_l419) && (inpThreshold <= CICC1851_when_SuperResolutionPart2_l428));
  assign when_SuperResolutionPart2_l430 = (inpThreshold <= CICC1851_when_SuperResolutionPart2_l419);
  assign when_SuperResolutionPart2_l431 = (inpThreshold <= CICC1851_when_SuperResolutionPart2_l419);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_valid = diffStage_controlPipe_fork_io_outputs_0_valid;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_payload_frameStart = diffStage_controlPipe_payload_frameStart;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_payload_rowEnd = diffStage_controlPipe_payload_rowEnd;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_payload_passMode = diffStage_controlPipe_payload_passMode;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_payload_passValid = diffStage_controlPipe_payload_passValid;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceMode = CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceMode;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceValid = CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceValid;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_payload_mainCompare = diffStage_controlPipe_payload_mainCompare;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_payload_counterCompare = diffStage_controlPipe_payload_counterCompare;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_payload_mainDiff = CICC1851_when_SuperResolutionPart2_l419;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_payload_counterDiff = CICC1851_when_SuperResolutionPart2_l428;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceCompValid = CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceCompValid;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceMode = CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceMode;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag = CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_payload_oddValid = diffStage_controlPipe_payload_oddValid;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_ready = (! diffStage_controlPipe_fork_io_outputs_0_translated_rValid);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_valid = (diffStage_controlPipe_fork_io_outputs_0_translated_valid || diffStage_controlPipe_fork_io_outputs_0_translated_rValid);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_frameStart = (diffStage_controlPipe_fork_io_outputs_0_translated_rValid ? diffStage_controlPipe_fork_io_outputs_0_translated_rData_frameStart : diffStage_controlPipe_fork_io_outputs_0_translated_payload_frameStart);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_rowEnd = (diffStage_controlPipe_fork_io_outputs_0_translated_rValid ? diffStage_controlPipe_fork_io_outputs_0_translated_rData_rowEnd : diffStage_controlPipe_fork_io_outputs_0_translated_payload_rowEnd);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_passMode = (diffStage_controlPipe_fork_io_outputs_0_translated_rValid ? diffStage_controlPipe_fork_io_outputs_0_translated_rData_passMode : diffStage_controlPipe_fork_io_outputs_0_translated_payload_passMode);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_passValid = (diffStage_controlPipe_fork_io_outputs_0_translated_rValid ? diffStage_controlPipe_fork_io_outputs_0_translated_rData_passValid : diffStage_controlPipe_fork_io_outputs_0_translated_payload_passValid);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_onceMode = (diffStage_controlPipe_fork_io_outputs_0_translated_rValid ? diffStage_controlPipe_fork_io_outputs_0_translated_rData_onceMode : diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceMode);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_onceValid = (diffStage_controlPipe_fork_io_outputs_0_translated_rValid ? diffStage_controlPipe_fork_io_outputs_0_translated_rData_onceValid : diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceValid);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_mainCompare = (diffStage_controlPipe_fork_io_outputs_0_translated_rValid ? diffStage_controlPipe_fork_io_outputs_0_translated_rData_mainCompare : diffStage_controlPipe_fork_io_outputs_0_translated_payload_mainCompare);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_counterCompare = (diffStage_controlPipe_fork_io_outputs_0_translated_rValid ? diffStage_controlPipe_fork_io_outputs_0_translated_rData_counterCompare : diffStage_controlPipe_fork_io_outputs_0_translated_payload_counterCompare);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_mainDiff = (diffStage_controlPipe_fork_io_outputs_0_translated_rValid ? diffStage_controlPipe_fork_io_outputs_0_translated_rData_mainDiff : diffStage_controlPipe_fork_io_outputs_0_translated_payload_mainDiff);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_counterDiff = (diffStage_controlPipe_fork_io_outputs_0_translated_rValid ? diffStage_controlPipe_fork_io_outputs_0_translated_rData_counterDiff : diffStage_controlPipe_fork_io_outputs_0_translated_payload_counterDiff);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_twiceCompValid = (diffStage_controlPipe_fork_io_outputs_0_translated_rValid ? diffStage_controlPipe_fork_io_outputs_0_translated_rData_twiceCompValid : diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceCompValid);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_twiceMode = (diffStage_controlPipe_fork_io_outputs_0_translated_rValid ? diffStage_controlPipe_fork_io_outputs_0_translated_rData_twiceMode : diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceMode);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_inpValidFlag = (diffStage_controlPipe_fork_io_outputs_0_translated_rValid ? diffStage_controlPipe_fork_io_outputs_0_translated_rData_inpValidFlag : diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_oddValid = (diffStage_controlPipe_fork_io_outputs_0_translated_rValid ? diffStage_controlPipe_fork_io_outputs_0_translated_rData_oddValid : diffStage_controlPipe_fork_io_outputs_0_translated_payload_oddValid);
  always @(*) begin
    diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_ready = resultStage_controlPipe_ready;
    if(when_Stream_l368_31) begin
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_31 = (! resultStage_controlPipe_valid);
  assign resultStage_controlPipe_valid = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rValid;
  assign resultStage_controlPipe_payload_frameStart = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_frameStart;
  assign resultStage_controlPipe_payload_rowEnd = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_rowEnd;
  assign resultStage_controlPipe_payload_passMode = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_passMode;
  assign resultStage_controlPipe_payload_passValid = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_passValid;
  assign resultStage_controlPipe_payload_onceMode = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_onceMode;
  assign resultStage_controlPipe_payload_onceValid = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_onceValid;
  assign resultStage_controlPipe_payload_mainCompare = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_mainCompare;
  assign resultStage_controlPipe_payload_counterCompare = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_counterCompare;
  assign resultStage_controlPipe_payload_mainDiff = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_mainDiff;
  assign resultStage_controlPipe_payload_counterDiff = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_counterDiff;
  assign resultStage_controlPipe_payload_twiceCompValid = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_twiceCompValid;
  assign resultStage_controlPipe_payload_twiceMode = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_twiceMode;
  assign resultStage_controlPipe_payload_inpValidFlag = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_inpValidFlag;
  assign resultStage_controlPipe_payload_oddValid = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_oddValid;
  assign resultStage_pixelStream_valid = diffStage_controlPipe_fork_io_outputs_1_valid;
  always @(*) begin
    resultStage_pixelStream_payload = 8'h0;
    if(diffStage_controlPipe_fork_io_outputs_1_payload_passValid) begin
      if(diffStage_controlPipe_fork_io_outputs_1_payload_passMode) begin
        resultStage_pixelStream_payload = diffStage_mainTwoPixelStream_payload;
      end else begin
        resultStage_pixelStream_payload = diffStage_mainOnePixelStream_payload;
      end
    end
    if(diffStage_controlPipe_fork_io_outputs_1_payload_oddValid) begin
      resultStage_pixelStream_payload = diffStage_oddRowPixelStream_payload;
    end
    if(diffStage_controlPipe_fork_io_outputs_1_payload_onceValid) begin
      case(diffStage_controlPipe_fork_io_outputs_1_payload_onceMode)
        3'b000 : begin
          if(when_SuperResolutionPart2_l451) begin
            resultStage_pixelStream_payload = 8'h0;
          end else begin
            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload[7:0];
          end
        end
        3'b001 : begin
          if(when_SuperResolutionPart2_l455) begin
            resultStage_pixelStream_payload = 8'h0;
          end else begin
            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_2[7:0];
          end
        end
        3'b010 : begin
          if(when_SuperResolutionPart2_l459) begin
            resultStage_pixelStream_payload = 8'h0;
          end else begin
            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_4[7:0];
          end
        end
        3'b011 : begin
          if(when_SuperResolutionPart2_l463) begin
            resultStage_pixelStream_payload = 8'h0;
          end else begin
            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_6[7:0];
          end
        end
        3'b100 : begin
          resultStage_pixelStream_payload = diffStage_mainOnePixelStream_payload;
        end
        3'b101 : begin
          resultStage_pixelStream_payload = diffStage_mainTwoPixelStream_payload;
        end
        default : begin
        end
      endcase
    end
    if(diffStage_controlPipe_fork_io_outputs_1_payload_twiceCompValid) begin
      case(diffStage_controlPipe_fork_io_outputs_1_payload_twiceMode)
        3'b000 : begin
          if(when_SuperResolutionPart2_l474) begin
            resultStage_pixelStream_payload = 8'h0;
          end else begin
            if(when_SuperResolutionPart2_l477) begin
              resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_8[7:0];
            end else begin
              resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_10[7:0];
            end
          end
        end
        3'b001 : begin
          if(when_SuperResolutionPart2_l482) begin
            resultStage_pixelStream_payload = 8'h0;
          end else begin
            if(when_SuperResolutionPart2_l485) begin
              resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_12[7:0];
            end else begin
              resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_14[7:0];
            end
          end
        end
        3'b010 : begin
          resultStage_pixelStream_payload = diffStage_mainTwoPixelStream_payload;
        end
        3'b011 : begin
          if(when_SuperResolutionPart2_l491) begin
            resultStage_pixelStream_payload = 8'h0;
          end else begin
            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_16[7:0];
          end
        end
        3'b100 : begin
          resultStage_pixelStream_payload = diffStage_mainOnePixelStream_payload;
        end
        3'b101 : begin
          if(when_SuperResolutionPart2_l496) begin
            resultStage_pixelStream_payload = 8'h0;
          end else begin
            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_18[7:0];
          end
        end
        default : begin
        end
      endcase
    end
  end

  assign when_SuperResolutionPart2_l451 = (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart2_l455 = (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart2_l459 = (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart2_l463 = (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart2_l474 = ((inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff) && (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff));
  assign when_SuperResolutionPart2_l477 = (diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart2_l482 = ((inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff) && (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff));
  assign when_SuperResolutionPart2_l485 = (diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart2_l491 = (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart2_l496 = (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign resultStage_pixelStream_ready = (! resultStage_pixelStream_rValid);
  assign resultStage_pixelStream_s2mPipe_valid = (resultStage_pixelStream_valid || resultStage_pixelStream_rValid);
  assign resultStage_pixelStream_s2mPipe_payload = (resultStage_pixelStream_rValid ? resultStage_pixelStream_rData : resultStage_pixelStream_payload);
  always @(*) begin
    resultStage_pixelStream_s2mPipe_ready = resultStage_resultStream_ready;
    if(when_Stream_l368_32) begin
      resultStage_pixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_32 = (! resultStage_resultStream_valid);
  assign resultStage_resultStream_valid = resultStage_pixelStream_s2mPipe_rValid;
  assign resultStage_resultStream_payload = resultStage_pixelStream_s2mPipe_rData;
  assign CICC1851_resultStage_mainOnePixelStream_ready_2 = (CICC1851_resultStage_mainOnePixelStream_ready && CICC1851_resultStage_mainOnePixelStream_ready_1);
  assign CICC1851_resultStage_mainOnePixelStream_ready = ((((((resultStage_resultStream_valid && resultStage_mainOnePixelStream_valid) && resultStage_counterOnePixelStream_valid) && resultStage_mainTwoPixelStream_valid) && resultStage_counterTwoPixelStream_valid) && resultStage_controlPipe_valid) && resultStage_oddRowPixelStream_valid);
  assign resultStage_resultStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_mainOnePixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_counterOnePixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_mainTwoPixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_counterTwoPixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_controlPipe_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_oddRowPixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign when_Stream_l438 = ((((! resultStage_controlPipe_payload_passValid) && (! resultStage_controlPipe_payload_onceValid)) && (! resultStage_controlPipe_payload_twiceCompValid)) && (! resultStage_controlPipe_payload_oddValid));
  always @(*) begin
    resultsJoin_valid = CICC1851_resultStage_mainOnePixelStream_ready;
    if(when_Stream_l438) begin
      resultsJoin_valid = 1'b0;
    end
  end

  always @(*) begin
    CICC1851_resultStage_mainOnePixelStream_ready_1 = resultsJoin_ready;
    if(when_Stream_l438) begin
      CICC1851_resultStage_mainOnePixelStream_ready_1 = 1'b1;
    end
  end

  assign pixelsStream_valid = resultsJoin_valid;
  assign resultsJoin_ready = pixelsStream_ready;
  assign pixelsStream_payload_pixel = resultStage_resultStream_payload;
  assign pixelsStream_payload_frameStart = resultStage_controlPipe_payload_frameStart;
  assign pixelsStream_payload_rowEnd = resultStage_controlPipe_payload_rowEnd;
  assign pixelsStream_payload_inpValid = resultStage_controlPipe_payload_inpValidFlag;
  assign pixelsStream_ready = (! pixelsStream_rValid);
  assign pixelsStream_s2mPipe_valid = (pixelsStream_valid || pixelsStream_rValid);
  assign pixelsStream_s2mPipe_payload_pixel = (pixelsStream_rValid ? pixelsStream_rData_pixel : pixelsStream_payload_pixel);
  assign pixelsStream_s2mPipe_payload_frameStart = (pixelsStream_rValid ? pixelsStream_rData_frameStart : pixelsStream_payload_frameStart);
  assign pixelsStream_s2mPipe_payload_rowEnd = (pixelsStream_rValid ? pixelsStream_rData_rowEnd : pixelsStream_payload_rowEnd);
  assign pixelsStream_s2mPipe_payload_inpValid = (pixelsStream_rValid ? pixelsStream_rData_inpValid : pixelsStream_payload_inpValid);
  always @(*) begin
    pixelsStream_s2mPipe_ready = pixelsStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_33) begin
      pixelsStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_33 = (! pixelsStream_s2mPipe_m2sPipe_valid);
  assign pixelsStream_s2mPipe_m2sPipe_valid = pixelsStream_s2mPipe_rValid;
  assign pixelsStream_s2mPipe_m2sPipe_payload_pixel = pixelsStream_s2mPipe_rData_pixel;
  assign pixelsStream_s2mPipe_m2sPipe_payload_frameStart = pixelsStream_s2mPipe_rData_frameStart;
  assign pixelsStream_s2mPipe_m2sPipe_payload_rowEnd = pixelsStream_s2mPipe_rData_rowEnd;
  assign pixelsStream_s2mPipe_m2sPipe_payload_inpValid = pixelsStream_s2mPipe_rData_inpValid;
  assign pixelsStream_s2mPipe_m2sPipe_ready = pixelsOut_ready;
  assign controlStateMachine_wantExit = 1'b0;
  always @(*) begin
    controlStateMachine_wantStart = 1'b0;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_7_HOLD : begin
      end
      controlStateMachine_enumDef_7_PASS : begin
      end
      controlStateMachine_enumDef_7_ONCE : begin
      end
      controlStateMachine_enumDef_7_TWICE : begin
      end
      default : begin
        controlStateMachine_wantStart = 1'b1;
      end
    endcase
  end

  assign controlStateMachine_wantKill = 1'b0;
  assign when_SuperResolutionPart2_l761 = (((currentState == 3'b010) || (currentState == 3'b011)) || (currentState == 3'b100));
  assign controlStream_fire_4 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart2_l763 = (controlStream_fire_4 && (CICC1851_when_SuperResolutionPart2_l763 == CICC1851_when_SuperResolutionPart2_l763_1));
  assign controlStream_fire_5 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart2_l764 = ((outReachRowEnd && (CICC1851_when_SuperResolutionPart2_l764 == CICC1851_when_SuperResolutionPart2_l764_1)) && controlStream_fire_5);
  assign controlStream_fire_6 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart2_l766 = (controlStream_fire_6 && outReachRowEnd);
  assign controlStream_fire_7 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart2_l783 = (CICC1851_when_SuperResolutionPart2_l783 == 12'h0);
  assign when_SuperResolutionPart2_l785 = (CICC1851_when_SuperResolutionPart2_l785 == 12'h001);
  assign when_SuperResolutionPart2_l787 = (CICC1851_when_SuperResolutionPart2_l787 == 12'h002);
  assign when_SuperResolutionPart2_l789 = (CICC1851_when_SuperResolutionPart2_l789 == 12'h003);
  assign when_SuperResolutionPart2_l793 = (CICC1851_when_SuperResolutionPart2_l793 == 12'h0);
  assign when_SuperResolutionPart2_l796 = (CICC1851_when_SuperResolutionPart2_l796 == 12'h001);
  assign when_SuperResolutionPart2_l799 = (CICC1851_when_SuperResolutionPart2_l799 == 12'h002);
  assign when_SuperResolutionPart2_l802 = (CICC1851_when_SuperResolutionPart2_l802 == 12'h003);
  always @(*) begin
    controlStateMachine_stateNext = controlStateMachine_stateReg;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_7_HOLD : begin
        if(zeroInFourOutRow) begin
          if(passPixels_fire_13) begin
            if(threeInFourOutPixelAddr) begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_7_ONCE;
            end else begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_7_PASS;
            end
          end
        end else begin
          if(twoInFourOutRow) begin
            if(passPixels_fire_14) begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_7_PASS;
            end
          end else begin
            if(threeInFourOutRow) begin
              if(passPixels_fire_15) begin
                if(threeInFourOutPixelAddr) begin
                  if(willHoldToTwice) begin
                    controlStateMachine_stateNext = controlStateMachine_enumDef_7_TWICE;
                  end
                end else begin
                  controlStateMachine_stateNext = controlStateMachine_enumDef_7_ONCE;
                end
              end
            end
          end
        end
      end
      controlStateMachine_enumDef_7_PASS : begin
        if(controlStream_fire_8) begin
          if(oneInFourOutPixelAddr) begin
            if(oneInFourOutRow) begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_7_PASS;
            end else begin
              if(twoInFourOutRow) begin
                if(when_SuperResolutionPart2_l573) begin
                  controlStateMachine_stateNext = controlStateMachine_enumDef_7_HOLD;
                end else begin
                  controlStateMachine_stateNext = controlStateMachine_enumDef_7_PASS;
                end
              end else begin
                if(when_SuperResolutionPart2_l578) begin
                  controlStateMachine_stateNext = controlStateMachine_enumDef_7_HOLD;
                end else begin
                  controlStateMachine_stateNext = controlStateMachine_enumDef_7_PASS;
                end
              end
            end
          end else begin
            if(twoInFourOutPixelAddr) begin
              if(oneInFourOutRow) begin
                controlStateMachine_stateNext = controlStateMachine_enumDef_7_ONCE;
              end else begin
                if(twoInFourOutRow) begin
                  controlStateMachine_stateNext = controlStateMachine_enumDef_7_ONCE;
                end else begin
                  if(when_SuperResolutionPart2_l590) begin
                    controlStateMachine_stateNext = controlStateMachine_enumDef_7_HOLD;
                  end else begin
                    controlStateMachine_stateNext = controlStateMachine_enumDef_7_ONCE;
                  end
                end
              end
            end else begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_7_PASS;
            end
          end
        end
      end
      controlStateMachine_enumDef_7_ONCE : begin
        if(controlStream_fire_10) begin
          if(zeroInFourOutRow) begin
            controlStateMachine_stateNext = controlStateMachine_enumDef_7_PASS;
          end else begin
            if(oneInFourOutRow) begin
              if(when_SuperResolutionPart2_l642) begin
                controlStateMachine_stateNext = controlStateMachine_enumDef_7_HOLD;
              end else begin
                controlStateMachine_stateNext = controlStateMachine_enumDef_7_PASS;
              end
            end else begin
              if(twoInFourOutRow) begin
                if(outReachRowEnd) begin
                  if(when_SuperResolutionPart2_l647) begin
                    controlStateMachine_stateNext = controlStateMachine_enumDef_7_HOLD;
                  end else begin
                    controlStateMachine_stateNext = controlStateMachine_enumDef_7_ONCE;
                  end
                end else begin
                  controlStateMachine_stateNext = controlStateMachine_enumDef_7_PASS;
                end
              end else begin
                if(twoInFourOutPixelAddr) begin
                  if(when_SuperResolutionPart2_l653) begin
                    controlStateMachine_stateNext = controlStateMachine_enumDef_7_HOLD;
                  end else begin
                    controlStateMachine_stateNext = controlStateMachine_enumDef_7_TWICE;
                  end
                end else begin
                  controlStateMachine_stateNext = controlStateMachine_enumDef_7_ONCE;
                end
              end
            end
          end
        end
      end
      controlStateMachine_enumDef_7_TWICE : begin
        if(controlStream_fire_11) begin
          if(outReachRowEnd) begin
            if(outReachFinalRow) begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_7_HOLD;
            end else begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_7_PASS;
            end
          end else begin
            controlStateMachine_stateNext = controlStateMachine_enumDef_7_ONCE;
          end
        end
      end
      default : begin
      end
    endcase
    if(controlStateMachine_wantStart) begin
      controlStateMachine_stateNext = controlStateMachine_enumDef_7_HOLD;
    end
    if(controlStateMachine_wantKill) begin
      controlStateMachine_stateNext = controlStateMachine_enumDef_7_BOOT;
    end
  end

  assign passPixels_fire_13 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_14 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_15 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_16 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart2_l560 = (CICC1851_when_SuperResolutionPart2_l560 == CICC1851_when_SuperResolutionPart2_l560_1);
  assign controlStream_fire_8 = (controlStream_valid && controlStream_ready);
  assign passPixels_fire_17 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart2_l573 = ((((oddBufferRow && (! holdBuffer)) && willPassToHoldCaseOne) && (! passPixels_fire_17)) && (! bufferReuse));
  assign passPixels_fire_18 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart2_l578 = (((((! oddBufferRow) && (! holdBuffer)) && willPassToHoldCaseOne) && (! passPixels_fire_18)) && (! bufferReuse));
  assign when_SuperResolutionPart2_l585 = ((oddBufferRow && (! holdBuffer)) && (! bufferReachRowEnd));
  assign when_SuperResolutionPart2_l588 = (((! oddBufferRow) && (! bufferReuse)) && (! bufferReachRowEnd));
  assign passPixels_fire_19 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart2_l590 = (((((! oddBufferRow) && (! holdBuffer)) && (! bufferReuse)) && (willPassToHoldCaseTwo || holdWillPassToHoldCaseTwo)) && (! passPixels_fire_19));
  assign when_SuperResolutionPart2_l602 = (poping && (CICC1851_when_SuperResolutionPart2_l602 == CICC1851_when_SuperResolutionPart2_l602_1));
  assign when_SuperResolutionPart2_l603 = (pushAndPoping && (CICC1851_when_SuperResolutionPart2_l603 == CICC1851_when_SuperResolutionPart2_l603_1));
  assign when_SuperResolutionPart2_l605 = (poping && (CICC1851_when_SuperResolutionPart2_l605 == CICC1851_when_SuperResolutionPart2_l605_1));
  assign when_SuperResolutionPart2_l606 = (pushAndPoping && (CICC1851_when_SuperResolutionPart2_l606 == CICC1851_when_SuperResolutionPart2_l606_1));
  assign when_SuperResolutionPart2_l609 = (CICC1851_when_SuperResolutionPart2_l609 == 12'h0);
  assign controlStream_fire_9 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart2_l630 = (frameStart && controlStream_fire_9);
  assign controlStream_fire_10 = (controlStream_valid && controlStream_ready);
  assign passPixels_fire_20 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart2_l642 = (((outReachRowEnd && willOnceToHoldCaseOne) && (bufferWAddr_value == 11'h0)) && (! passPixels_fire_20));
  assign passPixels_fire_21 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart2_l647 = (((bufferWAddr_value == 11'h0) && (! passPixels_fire_21)) && willOnceToHoldCaseTwo);
  assign passPixels_fire_22 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart2_l653 = ((((! oddBufferRow) && willOnceToHoldCaseThree) && (! passPixels_fire_22)) && (! bufferReuse));
  assign passPixels_fire_23 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart2_l662 = (passPixels_fire_23 && bufferReachRowEnd);
  assign when_SuperResolutionPart2_l667 = (poping && (CICC1851_when_SuperResolutionPart2_l667 == CICC1851_when_SuperResolutionPart2_l667_2));
  assign when_SuperResolutionPart2_l668 = (pushAndPoping && (CICC1851_when_SuperResolutionPart2_l668 == CICC1851_when_SuperResolutionPart2_l668_1));
  assign controlStream_fire_11 = (controlStream_valid && controlStream_ready);
  assign currentState = controlStateMachine_stateReg;
  always @(posedge clk or negedge resetn) begin
    if(!resetn) begin
      inpTwoDone <= 1'b0;
      readDone <= 1'b0;
      startRead <= 1'b0;
      slaveStart <= 1'b0;
      frameStart <= 1'b0;
      inpThreshold <= 8'h80;
      bmpWidth <= 10'h3c0;
      bmpHeight <= 10'h21c;
      holdBuffer <= 1'b0;
      writeDone <= 1'b0;
      bufferRowCount_value <= 11'h0;
      bufferReuse <= 1'b0;
      bufferEnable <= 1'b0;
      bufferSwitch <= 2'b00;
      nextRowBuffer <= 1'b1;
      bufferWAddr_value <= 11'h0;
      outPixelAddr_value <= 12'h0;
      outRowCount_value <= 12'h0;
      alreadySendRow_value <= 12'h0;
      alreadySendCountInRow_value <= 12'h0;
      alreadyReachRowEnd <= 1'b0;
      alreadyReachFinalRow <= 1'b0;
      outReachRowEnd <= 1'b0;
      outReachFinalRow <= 1'b0;
      bufferReachRowEnd <= 1'b0;
      bufferReachFinalRow <= 1'b0;
      oddBufferRow <= 1'b0;
      zeroInFourOutPixelAddr <= 1'b1;
      oneInFourOutPixelAddr <= 1'b0;
      twoInFourOutPixelAddr <= 1'b0;
      threeInFourOutPixelAddr <= 1'b0;
      zeroInFourOutRow <= 1'b1;
      oneInFourOutRow <= 1'b0;
      twoInFourOutRow <= 1'b0;
      threeInFourOutRow <= 1'b0;
      willHoldToTwice <= 1'b0;
      willPassToHoldCaseOne <= 1'b0;
      willPassToHoldCaseTwo <= 1'b0;
      holdWillPassToHoldCaseTwo <= 1'b0;
      willOnceToHoldCaseOne <= 1'b0;
      willOnceToHoldCaseTwo <= 1'b0;
      willOnceToHoldCaseThree <= 1'b0;
      pixelsIn_rValid <= 1'b0;
      pixelsIn_s2mPipe_rValid <= 1'b0;
      mainAddrOneStream_rValid <= 1'b0;
      mainAddrOneStream_s2mPipe_rValid <= 1'b0;
      CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_mainOnePixelStream_valid <= 1'b0;
      counterAddrOneStream_rValid <= 1'b0;
      counterAddrOneStream_s2mPipe_rValid <= 1'b0;
      CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_counterOnePixelStream_valid <= 1'b0;
      mainAddrTwoStream_rValid <= 1'b0;
      mainAddrTwoStream_s2mPipe_rValid <= 1'b0;
      CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_mainTwoPixelStream_valid <= 1'b0;
      counterAddrTwoStream_rValid <= 1'b0;
      counterAddrTwoStream_s2mPipe_rValid <= 1'b0;
      CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_counterTwoPixelStream_valid <= 1'b0;
      oddAddrStream_rValid <= 1'b0;
      oddAddrStream_s2mPipe_rValid <= 1'b0;
      CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_oddRowPixelStream_valid <= 1'b0;
      controlStream_rValid <= 1'b0;
      controlStream_s2mPipe_rValid <= 1'b0;
      controlStream_s2mPipe_m2sPipe_rValid <= 1'b0;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rValid <= 1'b0;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rValid <= 1'b0;
      readStage_mainOnePixelStream_rValid <= 1'b0;
      readStage_mainOnePixelStream_s2mPipe_rValid <= 1'b0;
      readStage_counterOnePixelStream_rValid <= 1'b0;
      readStage_counterOnePixelStream_s2mPipe_rValid <= 1'b0;
      readStage_mainTwoPixelStream_rValid <= 1'b0;
      readStage_mainTwoPixelStream_s2mPipe_rValid <= 1'b0;
      readStage_counterTwoPixelStream_rValid <= 1'b0;
      readStage_counterTwoPixelStream_s2mPipe_rValid <= 1'b0;
      readStage_oddRowPixelStream_rValid <= 1'b0;
      readStage_oddRowPixelStream_s2mPipe_rValid <= 1'b0;
      readStage_controlPipe_translated_rValid <= 1'b0;
      readStage_controlPipe_translated_s2mPipe_rValid <= 1'b0;
      compareStage_mainOnePixelStream_rValid <= 1'b0;
      compareStage_mainOnePixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_counterOnePixelStream_rValid <= 1'b0;
      compareStage_counterOnePixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_mainTwoPixelStream_rValid <= 1'b0;
      compareStage_mainTwoPixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_counterTwoPixelStream_rValid <= 1'b0;
      compareStage_counterTwoPixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_oddRowPixelStream_rValid <= 1'b0;
      compareStage_oddRowPixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_controlPipe_translated_rValid <= 1'b0;
      compareStage_controlPipe_translated_s2mPipe_rValid <= 1'b0;
      diffStage_mainOnePixelStream_rValid <= 1'b0;
      diffStage_mainOnePixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_counterOnePixelStream_rValid <= 1'b0;
      diffStage_counterOnePixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_mainTwoPixelStream_rValid <= 1'b0;
      diffStage_mainTwoPixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_counterTwoPixelStream_rValid <= 1'b0;
      diffStage_counterTwoPixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_oddRowPixelStream_rValid <= 1'b0;
      diffStage_oddRowPixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_controlPipe_fork_io_outputs_0_translated_rValid <= 1'b0;
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rValid <= 1'b0;
      resultStage_pixelStream_rValid <= 1'b0;
      resultStage_pixelStream_s2mPipe_rValid <= 1'b0;
      pixelsStream_rValid <= 1'b0;
      pixelsStream_s2mPipe_rValid <= 1'b0;
      controlStateMachine_stateReg <= controlStateMachine_enumDef_7_BOOT;
    end else begin
      if(when_SuperResolutionPart2_l40) begin
        inpTwoDone <= 1'b0;
      end
      if(when_SuperResolutionPart2_l43) begin
        readDone <= 1'b0;
      end
      if(when_SuperResolutionPart2_l46) begin
        startRead <= 1'b1;
      end
      if(when_SuperResolutionPart2_l46_1) begin
        startRead <= 1'b0;
      end
      if(when_SuperResolutionPart2_l49) begin
        slaveStart <= 1'b1;
      end
      if(when_SuperResolutionPart2_l49_1) begin
        slaveStart <= 1'b0;
      end
      inpThreshold <= thresholdIn;
      bmpWidth <= widthIn;
      bmpHeight <= heightIn;
      if(when_SuperResolutionPart2_l64) begin
        holdBuffer <= 1'b0;
      end
      if(when_SuperResolutionPart2_l67) begin
        writeDone <= 1'b0;
      end
      bufferRowCount_value <= bufferRowCount_valueNext;
      if(inpTwoDone) begin
        bufferReuse <= 1'b0;
      end
      if(when_SuperResolutionPart2_l76) begin
        bufferEnable <= 1'b1;
      end
      if(when_SuperResolutionPart2_l76_1) begin
        bufferEnable <= 1'b0;
      end
      if(when_SuperResolutionPart2_l82) begin
        nextRowBuffer <= 1'b1;
      end
      bufferWAddr_value <= bufferWAddr_valueNext;
      outPixelAddr_value <= outPixelAddr_valueNext;
      outRowCount_value <= outRowCount_valueNext;
      alreadySendRow_value <= alreadySendRow_valueNext;
      alreadySendCountInRow_value <= alreadySendCountInRow_valueNext;
      if(when_SuperResolutionPart2_l106) begin
        oddBufferRow <= 1'b0;
      end
      if(when_SuperResolutionPart2_l108) begin
        zeroInFourOutPixelAddr <= 1'b1;
      end
      if(when_SuperResolutionPart2_l109) begin
        oneInFourOutPixelAddr <= 1'b0;
      end
      if(when_SuperResolutionPart2_l110) begin
        twoInFourOutPixelAddr <= 1'b0;
      end
      if(when_SuperResolutionPart2_l111) begin
        threeInFourOutPixelAddr <= 1'b0;
      end
      if(when_SuperResolutionPart2_l113) begin
        zeroInFourOutRow <= 1'b1;
      end
      if(when_SuperResolutionPart2_l114) begin
        oneInFourOutRow <= 1'b0;
      end
      if(when_SuperResolutionPart2_l115) begin
        twoInFourOutRow <= 1'b0;
      end
      if(when_SuperResolutionPart2_l116) begin
        threeInFourOutRow <= 1'b0;
      end
      if(when_SuperResolutionPart2_l120) begin
        willHoldToTwice <= 1'b0;
      end
      if(when_SuperResolutionPart2_l121) begin
        willPassToHoldCaseOne <= 1'b0;
      end
      if(when_SuperResolutionPart2_l122) begin
        willPassToHoldCaseTwo <= 1'b0;
      end
      if(when_SuperResolutionPart2_l123) begin
        holdWillPassToHoldCaseTwo <= 1'b0;
      end
      if(when_SuperResolutionPart2_l124) begin
        willOnceToHoldCaseOne <= 1'b0;
      end
      if(when_SuperResolutionPart2_l125) begin
        willOnceToHoldCaseTwo <= 1'b0;
      end
      if(when_SuperResolutionPart2_l126) begin
        willOnceToHoldCaseThree <= 1'b0;
      end
      if(when_SuperResolutionPart2_l134) begin
        bufferSwitch <= 2'b00;
      end
      if(pixelsIn_valid) begin
        pixelsIn_rValid <= 1'b1;
      end
      if(pixelsIn_s2mPipe_ready) begin
        pixelsIn_rValid <= 1'b0;
      end
      if(pixelsIn_s2mPipe_ready) begin
        pixelsIn_s2mPipe_rValid <= pixelsIn_s2mPipe_valid;
      end
      if(when_SuperResolutionPart2_l181) begin
        bufferReachRowEnd <= 1'b1;
      end
      if(when_SuperResolutionPart2_l182) begin
        bufferReachFinalRow <= 1'b1;
      end
      if(when_SuperResolutionPart2_l185) begin
        if(bufferReachFinalRow) begin
          bufferReachRowEnd <= 1'b0;
          bufferReachFinalRow <= 1'b0;
          bufferReuse <= 1'b1;
        end else begin
          bufferReachRowEnd <= 1'b0;
        end
        if(when_SuperResolutionPart2_l195) begin
          oddBufferRow <= 1'b1;
        end else begin
          oddBufferRow <= 1'b0;
        end
      end
      if(when_SuperResolutionPart2_l200) begin
        if(when_SuperResolutionPart2_l201) begin
          bufferSwitch <= 2'b01;
        end else begin
          if(nextRowBuffer) begin
            bufferSwitch <= (bufferSwitch + 2'b01);
          end else begin
            bufferSwitch <= (bufferSwitch - 2'b01);
          end
        end
      end
      if(when_SuperResolutionPart2_l207) begin
        if(when_SuperResolutionPart2_l208) begin
          holdBuffer <= 1'b1;
          bufferEnable <= 1'b0;
        end
        if(when_SuperResolutionPart2_l212) begin
          writeDone <= 1'b1;
          bufferEnable <= 1'b0;
        end
      end
      if(when_SuperResolutionPart2_l218) begin
        holdBuffer <= 1'b0;
        if(when_SuperResolutionPart2_l220) begin
          nextRowBuffer <= (! nextRowBuffer);
        end
      end
      if(when_SuperResolutionPart2_l224) begin
        frameStart <= 1'b1;
      end
      if(when_SuperResolutionPart2_l234) begin
        alreadyReachRowEnd <= 1'b1;
      end
      if(when_SuperResolutionPart2_l235) begin
        alreadyReachFinalRow <= 1'b1;
      end
      if(pixelsOut_fire_2) begin
        if(alreadyReachRowEnd) begin
          alreadyReachRowEnd <= 1'b0;
          if(alreadyReachFinalRow) begin
            alreadyReachFinalRow <= 1'b0;
          end
        end
      end
      if(when_SuperResolutionPart2_l246) begin
        inpTwoDone <= 1'b1;
      end
      if(mainAddrOneStream_valid) begin
        mainAddrOneStream_rValid <= 1'b1;
      end
      if(mainAddrOneStream_s2mPipe_ready) begin
        mainAddrOneStream_rValid <= 1'b0;
      end
      if(mainAddrOneStream_s2mPipe_ready) begin
        mainAddrOneStream_s2mPipe_rValid <= mainAddrOneStream_s2mPipe_valid;
      end
      if(CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(mainAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_2 <= mainAddrOneStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_1) begin
        CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_1) begin
        CICC1851_readStage_mainOnePixelStream_valid <= (CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready || CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_3);
      end
      if(counterAddrOneStream_valid) begin
        counterAddrOneStream_rValid <= 1'b1;
      end
      if(counterAddrOneStream_s2mPipe_ready) begin
        counterAddrOneStream_rValid <= 1'b0;
      end
      if(counterAddrOneStream_s2mPipe_ready) begin
        counterAddrOneStream_s2mPipe_rValid <= counterAddrOneStream_s2mPipe_valid;
      end
      if(CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(counterAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_2 <= counterAddrOneStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_2) begin
        CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_2) begin
        CICC1851_readStage_counterOnePixelStream_valid <= (CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready || CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_3);
      end
      if(mainAddrTwoStream_valid) begin
        mainAddrTwoStream_rValid <= 1'b1;
      end
      if(mainAddrTwoStream_s2mPipe_ready) begin
        mainAddrTwoStream_rValid <= 1'b0;
      end
      if(mainAddrTwoStream_s2mPipe_ready) begin
        mainAddrTwoStream_s2mPipe_rValid <= mainAddrTwoStream_s2mPipe_valid;
      end
      if(CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(mainAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= mainAddrTwoStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_3) begin
        CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_3) begin
        CICC1851_readStage_mainTwoPixelStream_valid <= (CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready || CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_3);
      end
      if(counterAddrTwoStream_valid) begin
        counterAddrTwoStream_rValid <= 1'b1;
      end
      if(counterAddrTwoStream_s2mPipe_ready) begin
        counterAddrTwoStream_rValid <= 1'b0;
      end
      if(counterAddrTwoStream_s2mPipe_ready) begin
        counterAddrTwoStream_s2mPipe_rValid <= counterAddrTwoStream_s2mPipe_valid;
      end
      if(CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(counterAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= counterAddrTwoStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_4) begin
        CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_4) begin
        CICC1851_readStage_counterTwoPixelStream_valid <= (CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready || CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_3);
      end
      if(oddAddrStream_valid) begin
        oddAddrStream_rValid <= 1'b1;
      end
      if(oddAddrStream_s2mPipe_ready) begin
        oddAddrStream_rValid <= 1'b0;
      end
      if(oddAddrStream_s2mPipe_ready) begin
        oddAddrStream_s2mPipe_rValid <= oddAddrStream_s2mPipe_valid;
      end
      if(CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(oddAddrStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_2 <= oddAddrStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_5) begin
        CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_5) begin
        CICC1851_readStage_oddRowPixelStream_valid <= (CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready || CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_3);
      end
      if(controlStream_valid) begin
        controlStream_rValid <= 1'b1;
      end
      if(controlStream_s2mPipe_ready) begin
        controlStream_rValid <= 1'b0;
      end
      if(controlStream_s2mPipe_ready) begin
        controlStream_s2mPipe_rValid <= controlStream_s2mPipe_valid;
      end
      if(controlStream_s2mPipe_m2sPipe_ready) begin
        controlStream_s2mPipe_m2sPipe_rValid <= controlStream_s2mPipe_m2sPipe_valid;
      end
      if(controlStream_s2mPipe_m2sPipe_m2sPipe_valid) begin
        controlStream_s2mPipe_m2sPipe_m2sPipe_rValid <= 1'b1;
      end
      if(controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready) begin
        controlStream_s2mPipe_m2sPipe_m2sPipe_rValid <= 1'b0;
      end
      if(controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready) begin
        controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_valid;
      end
      if(readStage_mainOnePixelStream_valid) begin
        readStage_mainOnePixelStream_rValid <= 1'b1;
      end
      if(readStage_mainOnePixelStream_s2mPipe_ready) begin
        readStage_mainOnePixelStream_rValid <= 1'b0;
      end
      if(readStage_mainOnePixelStream_s2mPipe_ready) begin
        readStage_mainOnePixelStream_s2mPipe_rValid <= readStage_mainOnePixelStream_s2mPipe_valid;
      end
      if(readStage_counterOnePixelStream_valid) begin
        readStage_counterOnePixelStream_rValid <= 1'b1;
      end
      if(readStage_counterOnePixelStream_s2mPipe_ready) begin
        readStage_counterOnePixelStream_rValid <= 1'b0;
      end
      if(readStage_counterOnePixelStream_s2mPipe_ready) begin
        readStage_counterOnePixelStream_s2mPipe_rValid <= readStage_counterOnePixelStream_s2mPipe_valid;
      end
      if(readStage_mainTwoPixelStream_valid) begin
        readStage_mainTwoPixelStream_rValid <= 1'b1;
      end
      if(readStage_mainTwoPixelStream_s2mPipe_ready) begin
        readStage_mainTwoPixelStream_rValid <= 1'b0;
      end
      if(readStage_mainTwoPixelStream_s2mPipe_ready) begin
        readStage_mainTwoPixelStream_s2mPipe_rValid <= readStage_mainTwoPixelStream_s2mPipe_valid;
      end
      if(readStage_counterTwoPixelStream_valid) begin
        readStage_counterTwoPixelStream_rValid <= 1'b1;
      end
      if(readStage_counterTwoPixelStream_s2mPipe_ready) begin
        readStage_counterTwoPixelStream_rValid <= 1'b0;
      end
      if(readStage_counterTwoPixelStream_s2mPipe_ready) begin
        readStage_counterTwoPixelStream_s2mPipe_rValid <= readStage_counterTwoPixelStream_s2mPipe_valid;
      end
      if(readStage_oddRowPixelStream_valid) begin
        readStage_oddRowPixelStream_rValid <= 1'b1;
      end
      if(readStage_oddRowPixelStream_s2mPipe_ready) begin
        readStage_oddRowPixelStream_rValid <= 1'b0;
      end
      if(readStage_oddRowPixelStream_s2mPipe_ready) begin
        readStage_oddRowPixelStream_s2mPipe_rValid <= readStage_oddRowPixelStream_s2mPipe_valid;
      end
      if(readStage_controlPipe_translated_valid) begin
        readStage_controlPipe_translated_rValid <= 1'b1;
      end
      if(readStage_controlPipe_translated_s2mPipe_ready) begin
        readStage_controlPipe_translated_rValid <= 1'b0;
      end
      if(readStage_controlPipe_translated_s2mPipe_ready) begin
        readStage_controlPipe_translated_s2mPipe_rValid <= readStage_controlPipe_translated_s2mPipe_valid;
      end
      if(compareStage_mainOnePixelStream_valid) begin
        compareStage_mainOnePixelStream_rValid <= 1'b1;
      end
      if(compareStage_mainOnePixelStream_s2mPipe_ready) begin
        compareStage_mainOnePixelStream_rValid <= 1'b0;
      end
      if(compareStage_mainOnePixelStream_s2mPipe_ready) begin
        compareStage_mainOnePixelStream_s2mPipe_rValid <= compareStage_mainOnePixelStream_s2mPipe_valid;
      end
      if(compareStage_counterOnePixelStream_valid) begin
        compareStage_counterOnePixelStream_rValid <= 1'b1;
      end
      if(compareStage_counterOnePixelStream_s2mPipe_ready) begin
        compareStage_counterOnePixelStream_rValid <= 1'b0;
      end
      if(compareStage_counterOnePixelStream_s2mPipe_ready) begin
        compareStage_counterOnePixelStream_s2mPipe_rValid <= compareStage_counterOnePixelStream_s2mPipe_valid;
      end
      if(compareStage_mainTwoPixelStream_valid) begin
        compareStage_mainTwoPixelStream_rValid <= 1'b1;
      end
      if(compareStage_mainTwoPixelStream_s2mPipe_ready) begin
        compareStage_mainTwoPixelStream_rValid <= 1'b0;
      end
      if(compareStage_mainTwoPixelStream_s2mPipe_ready) begin
        compareStage_mainTwoPixelStream_s2mPipe_rValid <= compareStage_mainTwoPixelStream_s2mPipe_valid;
      end
      if(compareStage_counterTwoPixelStream_valid) begin
        compareStage_counterTwoPixelStream_rValid <= 1'b1;
      end
      if(compareStage_counterTwoPixelStream_s2mPipe_ready) begin
        compareStage_counterTwoPixelStream_rValid <= 1'b0;
      end
      if(compareStage_counterTwoPixelStream_s2mPipe_ready) begin
        compareStage_counterTwoPixelStream_s2mPipe_rValid <= compareStage_counterTwoPixelStream_s2mPipe_valid;
      end
      if(compareStage_oddRowPixelStream_valid) begin
        compareStage_oddRowPixelStream_rValid <= 1'b1;
      end
      if(compareStage_oddRowPixelStream_s2mPipe_ready) begin
        compareStage_oddRowPixelStream_rValid <= 1'b0;
      end
      if(compareStage_oddRowPixelStream_s2mPipe_ready) begin
        compareStage_oddRowPixelStream_s2mPipe_rValid <= compareStage_oddRowPixelStream_s2mPipe_valid;
      end
      if(compareStage_controlPipe_translated_valid) begin
        compareStage_controlPipe_translated_rValid <= 1'b1;
      end
      if(compareStage_controlPipe_translated_s2mPipe_ready) begin
        compareStage_controlPipe_translated_rValid <= 1'b0;
      end
      if(compareStage_controlPipe_translated_s2mPipe_ready) begin
        compareStage_controlPipe_translated_s2mPipe_rValid <= compareStage_controlPipe_translated_s2mPipe_valid;
      end
      if(diffStage_mainOnePixelStream_valid) begin
        diffStage_mainOnePixelStream_rValid <= 1'b1;
      end
      if(diffStage_mainOnePixelStream_s2mPipe_ready) begin
        diffStage_mainOnePixelStream_rValid <= 1'b0;
      end
      if(diffStage_mainOnePixelStream_s2mPipe_ready) begin
        diffStage_mainOnePixelStream_s2mPipe_rValid <= diffStage_mainOnePixelStream_s2mPipe_valid;
      end
      if(diffStage_counterOnePixelStream_valid) begin
        diffStage_counterOnePixelStream_rValid <= 1'b1;
      end
      if(diffStage_counterOnePixelStream_s2mPipe_ready) begin
        diffStage_counterOnePixelStream_rValid <= 1'b0;
      end
      if(diffStage_counterOnePixelStream_s2mPipe_ready) begin
        diffStage_counterOnePixelStream_s2mPipe_rValid <= diffStage_counterOnePixelStream_s2mPipe_valid;
      end
      if(diffStage_mainTwoPixelStream_valid) begin
        diffStage_mainTwoPixelStream_rValid <= 1'b1;
      end
      if(diffStage_mainTwoPixelStream_s2mPipe_ready) begin
        diffStage_mainTwoPixelStream_rValid <= 1'b0;
      end
      if(diffStage_mainTwoPixelStream_s2mPipe_ready) begin
        diffStage_mainTwoPixelStream_s2mPipe_rValid <= diffStage_mainTwoPixelStream_s2mPipe_valid;
      end
      if(diffStage_counterTwoPixelStream_valid) begin
        diffStage_counterTwoPixelStream_rValid <= 1'b1;
      end
      if(diffStage_counterTwoPixelStream_s2mPipe_ready) begin
        diffStage_counterTwoPixelStream_rValid <= 1'b0;
      end
      if(diffStage_counterTwoPixelStream_s2mPipe_ready) begin
        diffStage_counterTwoPixelStream_s2mPipe_rValid <= diffStage_counterTwoPixelStream_s2mPipe_valid;
      end
      if(diffStage_oddRowPixelStream_valid) begin
        diffStage_oddRowPixelStream_rValid <= 1'b1;
      end
      if(diffStage_oddRowPixelStream_s2mPipe_ready) begin
        diffStage_oddRowPixelStream_rValid <= 1'b0;
      end
      if(diffStage_oddRowPixelStream_s2mPipe_ready) begin
        diffStage_oddRowPixelStream_s2mPipe_rValid <= diffStage_oddRowPixelStream_s2mPipe_valid;
      end
      if(diffStage_controlPipe_fork_io_outputs_0_translated_valid) begin
        diffStage_controlPipe_fork_io_outputs_0_translated_rValid <= 1'b1;
      end
      if(diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_ready) begin
        diffStage_controlPipe_fork_io_outputs_0_translated_rValid <= 1'b0;
      end
      if(diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_ready) begin
        diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rValid <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_valid;
      end
      if(resultStage_pixelStream_valid) begin
        resultStage_pixelStream_rValid <= 1'b1;
      end
      if(resultStage_pixelStream_s2mPipe_ready) begin
        resultStage_pixelStream_rValid <= 1'b0;
      end
      if(resultStage_pixelStream_s2mPipe_ready) begin
        resultStage_pixelStream_s2mPipe_rValid <= resultStage_pixelStream_s2mPipe_valid;
      end
      if(pixelsStream_valid) begin
        pixelsStream_rValid <= 1'b1;
      end
      if(pixelsStream_s2mPipe_ready) begin
        pixelsStream_rValid <= 1'b0;
      end
      if(pixelsStream_s2mPipe_ready) begin
        pixelsStream_s2mPipe_rValid <= pixelsStream_s2mPipe_valid;
      end
      if(when_SuperResolutionPart2_l761) begin
        if(when_SuperResolutionPart2_l763) begin
          outReachRowEnd <= 1'b1;
        end
        if(when_SuperResolutionPart2_l764) begin
          outReachFinalRow <= 1'b1;
        end
        if(when_SuperResolutionPart2_l766) begin
          if(outReachFinalRow) begin
            startRead <= 1'b0;
            readDone <= 1'b1;
            outReachRowEnd <= 1'b0;
            outReachFinalRow <= 1'b0;
          end else begin
            outReachRowEnd <= 1'b0;
          end
        end
        if(controlStream_fire_7) begin
          if(outReachRowEnd) begin
            outReachRowEnd <= 1'b0;
            if(when_SuperResolutionPart2_l783) begin
              oneInFourOutRow <= 1'b1;
            end else begin
              oneInFourOutRow <= 1'b0;
            end
            if(when_SuperResolutionPart2_l785) begin
              twoInFourOutRow <= 1'b1;
            end else begin
              twoInFourOutRow <= 1'b0;
            end
            if(when_SuperResolutionPart2_l787) begin
              threeInFourOutRow <= 1'b1;
            end else begin
              threeInFourOutRow <= 1'b0;
            end
            if(when_SuperResolutionPart2_l789) begin
              zeroInFourOutRow <= 1'b1;
            end else begin
              zeroInFourOutRow <= 1'b0;
            end
          end
          if(when_SuperResolutionPart2_l793) begin
            oneInFourOutPixelAddr <= 1'b1;
          end
          if(oneInFourOutPixelAddr) begin
            oneInFourOutPixelAddr <= 1'b0;
          end
          if(when_SuperResolutionPart2_l796) begin
            twoInFourOutPixelAddr <= 1'b1;
          end
          if(twoInFourOutPixelAddr) begin
            twoInFourOutPixelAddr <= 1'b0;
          end
          if(when_SuperResolutionPart2_l799) begin
            threeInFourOutPixelAddr <= 1'b1;
          end
          if(threeInFourOutPixelAddr) begin
            threeInFourOutPixelAddr <= 1'b0;
          end
          if(when_SuperResolutionPart2_l802) begin
            zeroInFourOutPixelAddr <= 1'b1;
          end
          if(zeroInFourOutPixelAddr) begin
            zeroInFourOutPixelAddr <= 1'b0;
          end
        end
      end
      controlStateMachine_stateReg <= controlStateMachine_stateNext;
      case(controlStateMachine_stateReg)
        controlStateMachine_enumDef_7_HOLD : begin
          if(zeroInFourOutRow) begin
            if(passPixels_fire_13) begin
              if(!threeInFourOutPixelAddr) begin
                holdWillPassToHoldCaseTwo <= 1'b1;
              end
            end
          end else begin
            if(!twoInFourOutRow) begin
              if(threeInFourOutRow) begin
                if(passPixels_fire_15) begin
                  if(threeInFourOutPixelAddr) begin
                    if(willHoldToTwice) begin
                      willHoldToTwice <= 1'b0;
                    end
                  end
                end
              end
            end
          end
          if(passPixels_fire_16) begin
            if(when_SuperResolutionPart2_l560) begin
              willHoldToTwice <= 1'b1;
            end else begin
              willHoldToTwice <= 1'b0;
            end
          end
        end
        controlStateMachine_enumDef_7_PASS : begin
          if(controlStream_fire_8) begin
            if(!oneInFourOutPixelAddr) begin
              if(twoInFourOutPixelAddr) begin
                if(oneInFourOutRow) begin
                  if(when_SuperResolutionPart2_l585) begin
                    willOnceToHoldCaseOne <= 1'b1;
                  end
                end else begin
                  if(twoInFourOutRow) begin
                    if(when_SuperResolutionPart2_l588) begin
                      willOnceToHoldCaseTwo <= 1'b1;
                    end
                  end else begin
                    if(when_SuperResolutionPart2_l590) begin
                      holdWillPassToHoldCaseTwo <= 1'b0;
                    end
                  end
                end
              end
            end
            willPassToHoldCaseOne <= 1'b0;
            willPassToHoldCaseTwo <= 1'b0;
          end
          if(when_SuperResolutionPart2_l602) begin
            willPassToHoldCaseOne <= 1'b1;
          end
          if(when_SuperResolutionPart2_l603) begin
            willPassToHoldCaseOne <= 1'b1;
          end
          if(when_SuperResolutionPart2_l605) begin
            willPassToHoldCaseTwo <= 1'b1;
          end
          if(when_SuperResolutionPart2_l606) begin
            willPassToHoldCaseTwo <= 1'b1;
          end
          if(when_SuperResolutionPart2_l630) begin
            frameStart <= 1'b0;
          end
        end
        controlStateMachine_enumDef_7_ONCE : begin
          if(controlStream_fire_10) begin
            willOnceToHoldCaseOne <= 1'b0;
            willOnceToHoldCaseTwo <= 1'b0;
            willOnceToHoldCaseThree <= 1'b0;
          end
          if(when_SuperResolutionPart2_l662) begin
            willOnceToHoldCaseOne <= 1'b0;
            willOnceToHoldCaseTwo <= 1'b0;
          end
          if(when_SuperResolutionPart2_l667) begin
            willOnceToHoldCaseThree <= 1'b1;
          end
          if(when_SuperResolutionPart2_l668) begin
            willOnceToHoldCaseThree <= 1'b1;
          end
        end
        controlStateMachine_enumDef_7_TWICE : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(posedge clk) begin
    startIn_regNext <= startIn;
    startIn_regNext_1 <= startIn;
    startIn_regNext_2 <= startIn;
    startIn_regNext_3 <= startIn;
    startIn_regNext_4 <= startIn;
    startIn_regNext_5 <= startIn;
    startIn_regNext_6 <= startIn;
    startIn_regNext_7 <= startIn;
    startIn_regNext_8 <= startIn;
    startIn_regNext_9 <= startIn;
    startIn_regNext_10 <= startIn;
    startIn_regNext_11 <= startIn;
    startIn_regNext_12 <= startIn;
    startIn_regNext_13 <= startIn;
    startIn_regNext_14 <= startIn;
    startIn_regNext_15 <= startIn;
    startIn_regNext_16 <= startIn;
    if(pixelsIn_ready) begin
      pixelsIn_rData_pixel <= pixelsIn_payload_pixel;
      pixelsIn_rData_frameStart <= pixelsIn_payload_frameStart;
      pixelsIn_rData_rowEnd <= pixelsIn_payload_rowEnd;
    end
    if(pixelsIn_s2mPipe_ready) begin
      pixelsIn_s2mPipe_rData_pixel <= pixelsIn_s2mPipe_payload_pixel;
      pixelsIn_s2mPipe_rData_frameStart <= pixelsIn_s2mPipe_payload_frameStart;
      pixelsIn_s2mPipe_rData_rowEnd <= pixelsIn_s2mPipe_payload_rowEnd;
    end
    if(mainAddrOneStream_ready) begin
      mainAddrOneStream_rData <= mainAddrOneStream_payload;
    end
    if(mainAddrOneStream_s2mPipe_ready) begin
      mainAddrOneStream_s2mPipe_rData <= mainAddrOneStream_s2mPipe_payload;
    end
    if(CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_mainOnePixelStream_payload_1 <= CICC1851_readStage_mainOnePixelStream_payload;
    end
    if(CICC1851_1) begin
      CICC1851_readStage_mainOnePixelStream_payload_2 <= (CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_mainOnePixelStream_payload_1 : CICC1851_readStage_mainOnePixelStream_payload);
    end
    if(counterAddrOneStream_ready) begin
      counterAddrOneStream_rData <= counterAddrOneStream_payload;
    end
    if(counterAddrOneStream_s2mPipe_ready) begin
      counterAddrOneStream_s2mPipe_rData <= counterAddrOneStream_s2mPipe_payload;
    end
    if(CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_counterOnePixelStream_payload_1 <= CICC1851_readStage_counterOnePixelStream_payload;
    end
    if(CICC1851_2) begin
      CICC1851_readStage_counterOnePixelStream_payload_2 <= (CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_counterOnePixelStream_payload_1 : CICC1851_readStage_counterOnePixelStream_payload);
    end
    if(mainAddrTwoStream_ready) begin
      mainAddrTwoStream_rData <= mainAddrTwoStream_payload;
    end
    if(mainAddrTwoStream_s2mPipe_ready) begin
      mainAddrTwoStream_s2mPipe_rData <= mainAddrTwoStream_s2mPipe_payload;
    end
    if(CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_mainTwoPixelStream_payload_1 <= CICC1851_readStage_mainTwoPixelStream_payload;
    end
    if(CICC1851_3) begin
      CICC1851_readStage_mainTwoPixelStream_payload_2 <= (CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_mainTwoPixelStream_payload_1 : CICC1851_readStage_mainTwoPixelStream_payload);
    end
    if(counterAddrTwoStream_ready) begin
      counterAddrTwoStream_rData <= counterAddrTwoStream_payload;
    end
    if(counterAddrTwoStream_s2mPipe_ready) begin
      counterAddrTwoStream_s2mPipe_rData <= counterAddrTwoStream_s2mPipe_payload;
    end
    if(CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_counterTwoPixelStream_payload_1 <= CICC1851_readStage_counterTwoPixelStream_payload;
    end
    if(CICC1851_4) begin
      CICC1851_readStage_counterTwoPixelStream_payload_2 <= (CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_counterTwoPixelStream_payload_1 : CICC1851_readStage_counterTwoPixelStream_payload);
    end
    if(oddAddrStream_ready) begin
      oddAddrStream_rData <= oddAddrStream_payload;
    end
    if(oddAddrStream_s2mPipe_ready) begin
      oddAddrStream_s2mPipe_rData <= oddAddrStream_s2mPipe_payload;
    end
    if(CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_oddRowPixelStream_payload_1 <= CICC1851_readStage_oddRowPixelStream_payload;
    end
    if(CICC1851_5) begin
      CICC1851_readStage_oddRowPixelStream_payload_2 <= (CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_oddRowPixelStream_payload_1 : CICC1851_readStage_oddRowPixelStream_payload);
    end
    if(controlStream_ready) begin
      controlStream_rData_frameStart <= controlStream_payload_frameStart;
      controlStream_rData_rowEnd <= controlStream_payload_rowEnd;
      controlStream_rData_passMode <= controlStream_payload_passMode;
      controlStream_rData_passValid <= controlStream_payload_passValid;
      controlStream_rData_onceMode <= controlStream_payload_onceMode;
      controlStream_rData_onceValid <= controlStream_payload_onceValid;
      controlStream_rData_mainCompare <= controlStream_payload_mainCompare;
      controlStream_rData_counterCompare <= controlStream_payload_counterCompare;
      controlStream_rData_mainDiff <= controlStream_payload_mainDiff;
      controlStream_rData_counterDiff <= controlStream_payload_counterDiff;
      controlStream_rData_twiceCompValid <= controlStream_payload_twiceCompValid;
      controlStream_rData_twiceMode <= controlStream_payload_twiceMode;
      controlStream_rData_inpValidFlag <= controlStream_payload_inpValidFlag;
      controlStream_rData_oddValid <= controlStream_payload_oddValid;
    end
    if(controlStream_s2mPipe_ready) begin
      controlStream_s2mPipe_rData_frameStart <= controlStream_s2mPipe_payload_frameStart;
      controlStream_s2mPipe_rData_rowEnd <= controlStream_s2mPipe_payload_rowEnd;
      controlStream_s2mPipe_rData_passMode <= controlStream_s2mPipe_payload_passMode;
      controlStream_s2mPipe_rData_passValid <= controlStream_s2mPipe_payload_passValid;
      controlStream_s2mPipe_rData_onceMode <= controlStream_s2mPipe_payload_onceMode;
      controlStream_s2mPipe_rData_onceValid <= controlStream_s2mPipe_payload_onceValid;
      controlStream_s2mPipe_rData_mainCompare <= controlStream_s2mPipe_payload_mainCompare;
      controlStream_s2mPipe_rData_counterCompare <= controlStream_s2mPipe_payload_counterCompare;
      controlStream_s2mPipe_rData_mainDiff <= controlStream_s2mPipe_payload_mainDiff;
      controlStream_s2mPipe_rData_counterDiff <= controlStream_s2mPipe_payload_counterDiff;
      controlStream_s2mPipe_rData_twiceCompValid <= controlStream_s2mPipe_payload_twiceCompValid;
      controlStream_s2mPipe_rData_twiceMode <= controlStream_s2mPipe_payload_twiceMode;
      controlStream_s2mPipe_rData_inpValidFlag <= controlStream_s2mPipe_payload_inpValidFlag;
      controlStream_s2mPipe_rData_oddValid <= controlStream_s2mPipe_payload_oddValid;
    end
    if(controlStream_s2mPipe_m2sPipe_ready) begin
      controlStream_s2mPipe_m2sPipe_rData_frameStart <= controlStream_s2mPipe_m2sPipe_payload_frameStart;
      controlStream_s2mPipe_m2sPipe_rData_rowEnd <= controlStream_s2mPipe_m2sPipe_payload_rowEnd;
      controlStream_s2mPipe_m2sPipe_rData_passMode <= controlStream_s2mPipe_m2sPipe_payload_passMode;
      controlStream_s2mPipe_m2sPipe_rData_passValid <= controlStream_s2mPipe_m2sPipe_payload_passValid;
      controlStream_s2mPipe_m2sPipe_rData_onceMode <= controlStream_s2mPipe_m2sPipe_payload_onceMode;
      controlStream_s2mPipe_m2sPipe_rData_onceValid <= controlStream_s2mPipe_m2sPipe_payload_onceValid;
      controlStream_s2mPipe_m2sPipe_rData_mainCompare <= controlStream_s2mPipe_m2sPipe_payload_mainCompare;
      controlStream_s2mPipe_m2sPipe_rData_counterCompare <= controlStream_s2mPipe_m2sPipe_payload_counterCompare;
      controlStream_s2mPipe_m2sPipe_rData_mainDiff <= controlStream_s2mPipe_m2sPipe_payload_mainDiff;
      controlStream_s2mPipe_m2sPipe_rData_counterDiff <= controlStream_s2mPipe_m2sPipe_payload_counterDiff;
      controlStream_s2mPipe_m2sPipe_rData_twiceCompValid <= controlStream_s2mPipe_m2sPipe_payload_twiceCompValid;
      controlStream_s2mPipe_m2sPipe_rData_twiceMode <= controlStream_s2mPipe_m2sPipe_payload_twiceMode;
      controlStream_s2mPipe_m2sPipe_rData_inpValidFlag <= controlStream_s2mPipe_m2sPipe_payload_inpValidFlag;
      controlStream_s2mPipe_m2sPipe_rData_oddValid <= controlStream_s2mPipe_m2sPipe_payload_oddValid;
    end
    if(controlStream_s2mPipe_m2sPipe_m2sPipe_ready) begin
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_frameStart <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_frameStart;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_rowEnd <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_rowEnd;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_passMode <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passMode;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_passValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_onceMode <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceMode;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_onceValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_twiceCompValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceCompValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_twiceMode <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceMode;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_inpValidFlag <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_inpValidFlag;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_oddValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_oddValid;
    end
    if(controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready) begin
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_frameStart <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_frameStart;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_rowEnd <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_rowEnd;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_passMode <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_passMode;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_passValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_passValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_onceMode <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_onceMode;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_onceValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_onceValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_twiceCompValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_twiceCompValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_twiceMode <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_twiceMode;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_inpValidFlag <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_inpValidFlag;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_oddValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_oddValid;
    end
    if(readStage_mainOnePixelStream_ready) begin
      readStage_mainOnePixelStream_rData <= readStage_mainOnePixelStream_payload;
    end
    if(readStage_mainOnePixelStream_s2mPipe_ready) begin
      readStage_mainOnePixelStream_s2mPipe_rData <= readStage_mainOnePixelStream_s2mPipe_payload;
    end
    if(readStage_counterOnePixelStream_ready) begin
      readStage_counterOnePixelStream_rData <= readStage_counterOnePixelStream_payload;
    end
    if(readStage_counterOnePixelStream_s2mPipe_ready) begin
      readStage_counterOnePixelStream_s2mPipe_rData <= readStage_counterOnePixelStream_s2mPipe_payload;
    end
    if(readStage_mainTwoPixelStream_ready) begin
      readStage_mainTwoPixelStream_rData <= readStage_mainTwoPixelStream_payload;
    end
    if(readStage_mainTwoPixelStream_s2mPipe_ready) begin
      readStage_mainTwoPixelStream_s2mPipe_rData <= readStage_mainTwoPixelStream_s2mPipe_payload;
    end
    if(readStage_counterTwoPixelStream_ready) begin
      readStage_counterTwoPixelStream_rData <= readStage_counterTwoPixelStream_payload;
    end
    if(readStage_counterTwoPixelStream_s2mPipe_ready) begin
      readStage_counterTwoPixelStream_s2mPipe_rData <= readStage_counterTwoPixelStream_s2mPipe_payload;
    end
    if(readStage_oddRowPixelStream_ready) begin
      readStage_oddRowPixelStream_rData <= readStage_oddRowPixelStream_payload;
    end
    if(readStage_oddRowPixelStream_s2mPipe_ready) begin
      readStage_oddRowPixelStream_s2mPipe_rData <= readStage_oddRowPixelStream_s2mPipe_payload;
    end
    if(readStage_controlPipe_translated_ready) begin
      readStage_controlPipe_translated_rData_frameStart <= readStage_controlPipe_translated_payload_frameStart;
      readStage_controlPipe_translated_rData_rowEnd <= readStage_controlPipe_translated_payload_rowEnd;
      readStage_controlPipe_translated_rData_passMode <= readStage_controlPipe_translated_payload_passMode;
      readStage_controlPipe_translated_rData_passValid <= readStage_controlPipe_translated_payload_passValid;
      readStage_controlPipe_translated_rData_onceMode <= readStage_controlPipe_translated_payload_onceMode;
      readStage_controlPipe_translated_rData_onceValid <= readStage_controlPipe_translated_payload_onceValid;
      readStage_controlPipe_translated_rData_mainCompare <= readStage_controlPipe_translated_payload_mainCompare;
      readStage_controlPipe_translated_rData_counterCompare <= readStage_controlPipe_translated_payload_counterCompare;
      readStage_controlPipe_translated_rData_mainDiff <= readStage_controlPipe_translated_payload_mainDiff;
      readStage_controlPipe_translated_rData_counterDiff <= readStage_controlPipe_translated_payload_counterDiff;
      readStage_controlPipe_translated_rData_twiceCompValid <= readStage_controlPipe_translated_payload_twiceCompValid;
      readStage_controlPipe_translated_rData_twiceMode <= readStage_controlPipe_translated_payload_twiceMode;
      readStage_controlPipe_translated_rData_inpValidFlag <= readStage_controlPipe_translated_payload_inpValidFlag;
      readStage_controlPipe_translated_rData_oddValid <= readStage_controlPipe_translated_payload_oddValid;
    end
    if(readStage_controlPipe_translated_s2mPipe_ready) begin
      readStage_controlPipe_translated_s2mPipe_rData_frameStart <= readStage_controlPipe_translated_s2mPipe_payload_frameStart;
      readStage_controlPipe_translated_s2mPipe_rData_rowEnd <= readStage_controlPipe_translated_s2mPipe_payload_rowEnd;
      readStage_controlPipe_translated_s2mPipe_rData_passMode <= readStage_controlPipe_translated_s2mPipe_payload_passMode;
      readStage_controlPipe_translated_s2mPipe_rData_passValid <= readStage_controlPipe_translated_s2mPipe_payload_passValid;
      readStage_controlPipe_translated_s2mPipe_rData_onceMode <= readStage_controlPipe_translated_s2mPipe_payload_onceMode;
      readStage_controlPipe_translated_s2mPipe_rData_onceValid <= readStage_controlPipe_translated_s2mPipe_payload_onceValid;
      readStage_controlPipe_translated_s2mPipe_rData_mainCompare <= readStage_controlPipe_translated_s2mPipe_payload_mainCompare;
      readStage_controlPipe_translated_s2mPipe_rData_counterCompare <= readStage_controlPipe_translated_s2mPipe_payload_counterCompare;
      readStage_controlPipe_translated_s2mPipe_rData_mainDiff <= readStage_controlPipe_translated_s2mPipe_payload_mainDiff;
      readStage_controlPipe_translated_s2mPipe_rData_counterDiff <= readStage_controlPipe_translated_s2mPipe_payload_counterDiff;
      readStage_controlPipe_translated_s2mPipe_rData_twiceCompValid <= readStage_controlPipe_translated_s2mPipe_payload_twiceCompValid;
      readStage_controlPipe_translated_s2mPipe_rData_twiceMode <= readStage_controlPipe_translated_s2mPipe_payload_twiceMode;
      readStage_controlPipe_translated_s2mPipe_rData_inpValidFlag <= readStage_controlPipe_translated_s2mPipe_payload_inpValidFlag;
      readStage_controlPipe_translated_s2mPipe_rData_oddValid <= readStage_controlPipe_translated_s2mPipe_payload_oddValid;
    end
    if(compareStage_mainOnePixelStream_ready) begin
      compareStage_mainOnePixelStream_rData <= compareStage_mainOnePixelStream_payload;
    end
    if(compareStage_mainOnePixelStream_s2mPipe_ready) begin
      compareStage_mainOnePixelStream_s2mPipe_rData <= compareStage_mainOnePixelStream_s2mPipe_payload;
    end
    if(compareStage_counterOnePixelStream_ready) begin
      compareStage_counterOnePixelStream_rData <= compareStage_counterOnePixelStream_payload;
    end
    if(compareStage_counterOnePixelStream_s2mPipe_ready) begin
      compareStage_counterOnePixelStream_s2mPipe_rData <= compareStage_counterOnePixelStream_s2mPipe_payload;
    end
    if(compareStage_mainTwoPixelStream_ready) begin
      compareStage_mainTwoPixelStream_rData <= compareStage_mainTwoPixelStream_payload;
    end
    if(compareStage_mainTwoPixelStream_s2mPipe_ready) begin
      compareStage_mainTwoPixelStream_s2mPipe_rData <= compareStage_mainTwoPixelStream_s2mPipe_payload;
    end
    if(compareStage_counterTwoPixelStream_ready) begin
      compareStage_counterTwoPixelStream_rData <= compareStage_counterTwoPixelStream_payload;
    end
    if(compareStage_counterTwoPixelStream_s2mPipe_ready) begin
      compareStage_counterTwoPixelStream_s2mPipe_rData <= compareStage_counterTwoPixelStream_s2mPipe_payload;
    end
    if(compareStage_oddRowPixelStream_ready) begin
      compareStage_oddRowPixelStream_rData <= compareStage_oddRowPixelStream_payload;
    end
    if(compareStage_oddRowPixelStream_s2mPipe_ready) begin
      compareStage_oddRowPixelStream_s2mPipe_rData <= compareStage_oddRowPixelStream_s2mPipe_payload;
    end
    if(compareStage_controlPipe_translated_ready) begin
      compareStage_controlPipe_translated_rData_frameStart <= compareStage_controlPipe_translated_payload_frameStart;
      compareStage_controlPipe_translated_rData_rowEnd <= compareStage_controlPipe_translated_payload_rowEnd;
      compareStage_controlPipe_translated_rData_passMode <= compareStage_controlPipe_translated_payload_passMode;
      compareStage_controlPipe_translated_rData_passValid <= compareStage_controlPipe_translated_payload_passValid;
      compareStage_controlPipe_translated_rData_onceMode <= compareStage_controlPipe_translated_payload_onceMode;
      compareStage_controlPipe_translated_rData_onceValid <= compareStage_controlPipe_translated_payload_onceValid;
      compareStage_controlPipe_translated_rData_mainCompare <= compareStage_controlPipe_translated_payload_mainCompare;
      compareStage_controlPipe_translated_rData_counterCompare <= compareStage_controlPipe_translated_payload_counterCompare;
      compareStage_controlPipe_translated_rData_mainDiff <= compareStage_controlPipe_translated_payload_mainDiff;
      compareStage_controlPipe_translated_rData_counterDiff <= compareStage_controlPipe_translated_payload_counterDiff;
      compareStage_controlPipe_translated_rData_twiceCompValid <= compareStage_controlPipe_translated_payload_twiceCompValid;
      compareStage_controlPipe_translated_rData_twiceMode <= compareStage_controlPipe_translated_payload_twiceMode;
      compareStage_controlPipe_translated_rData_inpValidFlag <= compareStage_controlPipe_translated_payload_inpValidFlag;
      compareStage_controlPipe_translated_rData_oddValid <= compareStage_controlPipe_translated_payload_oddValid;
    end
    if(compareStage_controlPipe_translated_s2mPipe_ready) begin
      compareStage_controlPipe_translated_s2mPipe_rData_frameStart <= compareStage_controlPipe_translated_s2mPipe_payload_frameStart;
      compareStage_controlPipe_translated_s2mPipe_rData_rowEnd <= compareStage_controlPipe_translated_s2mPipe_payload_rowEnd;
      compareStage_controlPipe_translated_s2mPipe_rData_passMode <= compareStage_controlPipe_translated_s2mPipe_payload_passMode;
      compareStage_controlPipe_translated_s2mPipe_rData_passValid <= compareStage_controlPipe_translated_s2mPipe_payload_passValid;
      compareStage_controlPipe_translated_s2mPipe_rData_onceMode <= compareStage_controlPipe_translated_s2mPipe_payload_onceMode;
      compareStage_controlPipe_translated_s2mPipe_rData_onceValid <= compareStage_controlPipe_translated_s2mPipe_payload_onceValid;
      compareStage_controlPipe_translated_s2mPipe_rData_mainCompare <= compareStage_controlPipe_translated_s2mPipe_payload_mainCompare;
      compareStage_controlPipe_translated_s2mPipe_rData_counterCompare <= compareStage_controlPipe_translated_s2mPipe_payload_counterCompare;
      compareStage_controlPipe_translated_s2mPipe_rData_mainDiff <= compareStage_controlPipe_translated_s2mPipe_payload_mainDiff;
      compareStage_controlPipe_translated_s2mPipe_rData_counterDiff <= compareStage_controlPipe_translated_s2mPipe_payload_counterDiff;
      compareStage_controlPipe_translated_s2mPipe_rData_twiceCompValid <= compareStage_controlPipe_translated_s2mPipe_payload_twiceCompValid;
      compareStage_controlPipe_translated_s2mPipe_rData_twiceMode <= compareStage_controlPipe_translated_s2mPipe_payload_twiceMode;
      compareStage_controlPipe_translated_s2mPipe_rData_inpValidFlag <= compareStage_controlPipe_translated_s2mPipe_payload_inpValidFlag;
      compareStage_controlPipe_translated_s2mPipe_rData_oddValid <= compareStage_controlPipe_translated_s2mPipe_payload_oddValid;
    end
    if(diffStage_mainOnePixelStream_ready) begin
      diffStage_mainOnePixelStream_rData <= diffStage_mainOnePixelStream_payload;
    end
    if(diffStage_mainOnePixelStream_s2mPipe_ready) begin
      diffStage_mainOnePixelStream_s2mPipe_rData <= diffStage_mainOnePixelStream_s2mPipe_payload;
    end
    if(diffStage_counterOnePixelStream_ready) begin
      diffStage_counterOnePixelStream_rData <= diffStage_counterOnePixelStream_payload;
    end
    if(diffStage_counterOnePixelStream_s2mPipe_ready) begin
      diffStage_counterOnePixelStream_s2mPipe_rData <= diffStage_counterOnePixelStream_s2mPipe_payload;
    end
    if(diffStage_mainTwoPixelStream_ready) begin
      diffStage_mainTwoPixelStream_rData <= diffStage_mainTwoPixelStream_payload;
    end
    if(diffStage_mainTwoPixelStream_s2mPipe_ready) begin
      diffStage_mainTwoPixelStream_s2mPipe_rData <= diffStage_mainTwoPixelStream_s2mPipe_payload;
    end
    if(diffStage_counterTwoPixelStream_ready) begin
      diffStage_counterTwoPixelStream_rData <= diffStage_counterTwoPixelStream_payload;
    end
    if(diffStage_counterTwoPixelStream_s2mPipe_ready) begin
      diffStage_counterTwoPixelStream_s2mPipe_rData <= diffStage_counterTwoPixelStream_s2mPipe_payload;
    end
    if(diffStage_oddRowPixelStream_ready) begin
      diffStage_oddRowPixelStream_rData <= diffStage_oddRowPixelStream_payload;
    end
    if(diffStage_oddRowPixelStream_s2mPipe_ready) begin
      diffStage_oddRowPixelStream_s2mPipe_rData <= diffStage_oddRowPixelStream_s2mPipe_payload;
    end
    if(diffStage_controlPipe_fork_io_outputs_0_translated_ready) begin
      diffStage_controlPipe_fork_io_outputs_0_translated_rData_frameStart <= diffStage_controlPipe_fork_io_outputs_0_translated_payload_frameStart;
      diffStage_controlPipe_fork_io_outputs_0_translated_rData_rowEnd <= diffStage_controlPipe_fork_io_outputs_0_translated_payload_rowEnd;
      diffStage_controlPipe_fork_io_outputs_0_translated_rData_passMode <= diffStage_controlPipe_fork_io_outputs_0_translated_payload_passMode;
      diffStage_controlPipe_fork_io_outputs_0_translated_rData_passValid <= diffStage_controlPipe_fork_io_outputs_0_translated_payload_passValid;
      diffStage_controlPipe_fork_io_outputs_0_translated_rData_onceMode <= diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceMode;
      diffStage_controlPipe_fork_io_outputs_0_translated_rData_onceValid <= diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceValid;
      diffStage_controlPipe_fork_io_outputs_0_translated_rData_mainCompare <= diffStage_controlPipe_fork_io_outputs_0_translated_payload_mainCompare;
      diffStage_controlPipe_fork_io_outputs_0_translated_rData_counterCompare <= diffStage_controlPipe_fork_io_outputs_0_translated_payload_counterCompare;
      diffStage_controlPipe_fork_io_outputs_0_translated_rData_mainDiff <= diffStage_controlPipe_fork_io_outputs_0_translated_payload_mainDiff;
      diffStage_controlPipe_fork_io_outputs_0_translated_rData_counterDiff <= diffStage_controlPipe_fork_io_outputs_0_translated_payload_counterDiff;
      diffStage_controlPipe_fork_io_outputs_0_translated_rData_twiceCompValid <= diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceCompValid;
      diffStage_controlPipe_fork_io_outputs_0_translated_rData_twiceMode <= diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceMode;
      diffStage_controlPipe_fork_io_outputs_0_translated_rData_inpValidFlag <= diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag;
      diffStage_controlPipe_fork_io_outputs_0_translated_rData_oddValid <= diffStage_controlPipe_fork_io_outputs_0_translated_payload_oddValid;
    end
    if(diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_ready) begin
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_frameStart <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_frameStart;
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_rowEnd <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_rowEnd;
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_passMode <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_passMode;
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_passValid <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_passValid;
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_onceMode <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_onceMode;
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_onceValid <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_onceValid;
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_mainCompare <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_mainCompare;
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_counterCompare <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_counterCompare;
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_mainDiff <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_mainDiff;
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_counterDiff <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_counterDiff;
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_twiceCompValid <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_twiceCompValid;
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_twiceMode <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_twiceMode;
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_inpValidFlag <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_inpValidFlag;
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_oddValid <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_oddValid;
    end
    if(resultStage_pixelStream_ready) begin
      resultStage_pixelStream_rData <= resultStage_pixelStream_payload;
    end
    if(resultStage_pixelStream_s2mPipe_ready) begin
      resultStage_pixelStream_s2mPipe_rData <= resultStage_pixelStream_s2mPipe_payload;
    end
    if(pixelsStream_ready) begin
      pixelsStream_rData_pixel <= pixelsStream_payload_pixel;
      pixelsStream_rData_frameStart <= pixelsStream_payload_frameStart;
      pixelsStream_rData_rowEnd <= pixelsStream_payload_rowEnd;
      pixelsStream_rData_inpValid <= pixelsStream_payload_inpValid;
    end
    if(pixelsStream_s2mPipe_ready) begin
      pixelsStream_s2mPipe_rData_pixel <= pixelsStream_s2mPipe_payload_pixel;
      pixelsStream_s2mPipe_rData_frameStart <= pixelsStream_s2mPipe_payload_frameStart;
      pixelsStream_s2mPipe_rData_rowEnd <= pixelsStream_s2mPipe_payload_rowEnd;
      pixelsStream_s2mPipe_rData_inpValid <= pixelsStream_s2mPipe_payload_inpValid;
    end
  end


endmodule

module SuperResolutionPart1_2 (
  input               pixelsIn_valid,
  output reg          pixelsIn_ready,
  input      [7:0]    pixelsIn_payload_pixel,
  input               pixelsIn_payload_frameStart,
  input               pixelsIn_payload_rowEnd,
  input               startIn,
  input               inpTwoDoneIn,
  input               inpThreeDoneIn,
  output reg          pixelsOut_valid,
  input               pixelsOut_ready,
  output reg [7:0]    pixelsOut_payload_pixel,
  output reg          pixelsOut_payload_frameStart,
  output reg          pixelsOut_payload_rowEnd,
  output reg          startOut,
  output reg          inpDoneOut,
  input      [7:0]    thresholdIn,
  input      [9:0]    widthIn,
  input      [9:0]    heightIn,
  input               clk,
  input               resetn
);
  localparam controlStateMachine_enumDef_6_BOOT = 3'd0;
  localparam controlStateMachine_enumDef_6_HOLD = 3'd1;
  localparam controlStateMachine_enumDef_6_PASS = 3'd2;
  localparam controlStateMachine_enumDef_6_ONCE = 3'd3;
  localparam controlStateMachine_enumDef_6_TWICE = 3'd4;

  wire                diffStage_controlPipe_fork_io_outputs_0_ready;
  reg        [7:0]    CICC1851_lineBufferOne_port0;
  reg        [7:0]    CICC1851_lineBufferOne_port1;
  reg        [7:0]    CICC1851_lineBufferTwo_port0;
  reg        [7:0]    CICC1851_lineBufferTwo_port1;
  wire                diffStage_controlPipe_fork_io_input_ready;
  wire                diffStage_controlPipe_fork_io_outputs_0_valid;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_frameStart;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_rowEnd;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_passMode;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_passValid;
  wire       [2:0]    diffStage_controlPipe_fork_io_outputs_0_payload_onceMode;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_onceValid;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_mainCompare;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_counterCompare;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_payload_mainDiff;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_payload_counterDiff;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_twiceCompValid;
  wire       [2:0]    diffStage_controlPipe_fork_io_outputs_0_payload_twiceMode;
  wire                diffStage_controlPipe_fork_io_outputs_1_valid;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_frameStart;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_rowEnd;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_passMode;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_passValid;
  wire       [2:0]    diffStage_controlPipe_fork_io_outputs_1_payload_onceMode;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_onceValid;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_mainCompare;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_counterCompare;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_twiceCompValid;
  wire       [2:0]    diffStage_controlPipe_fork_io_outputs_1_payload_twiceMode;
  wire       [9:0]    CICC1851_bufferRowCount_valueNext;
  wire       [0:0]    CICC1851_bufferRowCount_valueNext_1;
  wire       [9:0]    CICC1851_bufferWAddr_valueNext;
  wire       [0:0]    CICC1851_bufferWAddr_valueNext_1;
  wire       [10:0]   CICC1851_outPixelAddr_valueNext;
  wire       [0:0]    CICC1851_outPixelAddr_valueNext_1;
  wire       [10:0]   CICC1851_outRowCount_valueNext;
  wire       [0:0]    CICC1851_outRowCount_valueNext_1;
  wire       [10:0]   CICC1851_mainAddrOne;
  wire       [10:0]   CICC1851_counterAddrOne;
  wire       [10:0]   CICC1851_mainAddrTwo;
  wire       [10:0]   CICC1851_counterAddrTwo;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_1;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_2;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_3;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_4;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_5;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_6;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_7;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_8;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_9;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_10;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_11;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_12;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_13;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_14;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_15;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_16;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_17;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_18;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_19;
  wire       [9:0]    CICC1851_when_SuperResolutionPart1_l421;
  wire       [9:0]    CICC1851_when_SuperResolutionPart1_l422;
  wire       [10:0]   CICC1851_when_SuperResolutionPart1_l447;
  wire       [7:0]    CICC1851_lineBufferTwo_port;
  wire                CICC1851_lineBufferTwo_port_1;
  wire       [7:0]    CICC1851_lineBufferOne_port;
  wire                CICC1851_lineBufferOne_port_1;
  wire       [10:0]   CICC1851_when_SuperResolutionPart1_l482;
  wire       [10:0]   CICC1851_when_SuperResolutionPart1_l484;
  wire       [10:0]   CICC1851_when_SuperResolutionPart1_l489;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l498;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l498_1;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l500;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l500_1;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l500_2;
  wire       [2:0]    CICC1851_when_SuperResolutionPart1_l500_3;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l510;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l510_1;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l510_2;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l511;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l511_1;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l511_2;
  wire       [10:0]   CICC1851_when_SuperResolutionPart1_l537;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l542;
  wire       [10:0]   CICC1851_when_SuperResolutionPart1_l542_1;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l542_2;
  wire       [10:0]   CICC1851_mainAddrOne_1;
  wire       [10:0]   CICC1851_mainAddrOne_2;
  wire       [10:0]   CICC1851_counterAddrOne_1;
  wire       [10:0]   CICC1851_counterAddrOne_2;
  wire       [11:0]   CICC1851_counterAddrOne_3;
  wire       [11:0]   CICC1851_counterAddrOne_4;
  wire       [11:0]   CICC1851_counterAddrOne_5;
  wire       [1:0]    CICC1851_counterAddrOne_6;
  wire       [0:0]    CICC1851_controls_onceMode;
  wire       [10:0]   CICC1851_mainAddrTwo_1;
  wire       [10:0]   CICC1851_mainAddrTwo_2;
  wire       [10:0]   CICC1851_counterAddrTwo_1;
  wire       [10:0]   CICC1851_counterAddrTwo_2;
  wire       [11:0]   CICC1851_counterAddrTwo_3;
  wire       [11:0]   CICC1851_counterAddrTwo_4;
  wire       [11:0]   CICC1851_counterAddrTwo_5;
  wire       [1:0]    CICC1851_counterAddrTwo_6;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l563;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l563_1;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l563_2;
  wire       [2:0]    CICC1851_when_SuperResolutionPart1_l563_3;
  wire       [1:0]    CICC1851_controls_onceMode_1;
  wire       [1:0]    CICC1851_controls_onceMode_2;
  wire       [10:0]   CICC1851_mainAddrOne_3;
  wire       [10:0]   CICC1851_mainAddrTwo_3;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l578;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l578_1;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l578_2;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l579;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l579_1;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l579_2;
  wire       [10:0]   CICC1851_mainAddrOne_4;
  wire       [10:0]   CICC1851_mainAddrOne_5;
  wire       [10:0]   CICC1851_mainAddrOne_6;
  wire       [10:0]   CICC1851_mainAddrOne_7;
  wire       [11:0]   CICC1851_counterAddrOne_7;
  wire       [11:0]   CICC1851_counterAddrOne_8;
  wire       [11:0]   CICC1851_counterAddrOne_9;
  wire       [1:0]    CICC1851_counterAddrOne_10;
  wire       [10:0]   CICC1851_mainAddrTwo_4;
  wire       [10:0]   CICC1851_mainAddrTwo_5;
  wire       [10:0]   CICC1851_mainAddrTwo_6;
  wire       [10:0]   CICC1851_mainAddrTwo_7;
  wire       [11:0]   CICC1851_counterAddrTwo_7;
  wire       [11:0]   CICC1851_counterAddrTwo_8;
  wire       [11:0]   CICC1851_counterAddrTwo_9;
  wire       [1:0]    CICC1851_counterAddrTwo_10;
  wire       [10:0]   CICC1851_mainAddrOne_8;
  wire       [10:0]   CICC1851_mainAddrOne_9;
  wire       [10:0]   CICC1851_counterAddrTwo_11;
  wire       [10:0]   CICC1851_counterAddrTwo_12;
  wire       [10:0]   CICC1851_mainAddrTwo_8;
  wire       [10:0]   CICC1851_mainAddrTwo_9;
  wire       [10:0]   CICC1851_counterAddrOne_11;
  wire       [10:0]   CICC1851_counterAddrOne_12;
  wire       [11:0]   CICC1851_mainAddrTwo_10;
  wire       [11:0]   CICC1851_mainAddrTwo_11;
  wire       [11:0]   CICC1851_mainAddrTwo_12;
  wire       [1:0]    CICC1851_mainAddrTwo_13;
  wire       [11:0]   CICC1851_counterAddrOne_13;
  wire       [11:0]   CICC1851_counterAddrOne_14;
  wire       [11:0]   CICC1851_counterAddrOne_15;
  wire       [1:0]    CICC1851_counterAddrOne_16;
  wire       [10:0]   CICC1851_mainAddrTwo_14;
  wire       [10:0]   CICC1851_mainAddrTwo_15;
  wire       [10:0]   CICC1851_counterAddrOne_17;
  wire       [10:0]   CICC1851_counterAddrOne_18;
  wire       [10:0]   CICC1851_mainAddrOne_10;
  wire       [10:0]   CICC1851_mainAddrOne_11;
  wire       [10:0]   CICC1851_counterAddrTwo_13;
  wire       [10:0]   CICC1851_counterAddrTwo_14;
  wire       [11:0]   CICC1851_mainAddrOne_12;
  wire       [11:0]   CICC1851_mainAddrOne_13;
  wire       [11:0]   CICC1851_mainAddrOne_14;
  wire       [1:0]    CICC1851_mainAddrOne_15;
  wire       [11:0]   CICC1851_counterAddrTwo_15;
  wire       [11:0]   CICC1851_counterAddrTwo_16;
  wire       [11:0]   CICC1851_counterAddrTwo_17;
  wire       [1:0]    CICC1851_counterAddrTwo_18;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l664;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l664_1;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l664_2;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l665;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l665_1;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l665_2;
  reg                 inpDone;
  wire                when_SuperResolutionPart1_l79;
  reg                 startIn_regNext;
  wire                when_SuperResolutionPart1_l79_1;
  reg                 readDone;
  wire                when_SuperResolutionPart1_l82;
  reg                 startRead;
  wire                when_SuperResolutionPart1_l85;
  wire                when_SuperResolutionPart1_l85_1;
  reg                 slaveStart;
  wire                pixelsIn_fire;
  wire                when_SuperResolutionPart1_l88;
  wire                when_SuperResolutionPart1_l88_1;
  reg                 frameStart;
  reg        [7:0]    inpThreshold;
  reg        [9:0]    bmpWidth;
  reg        [9:0]    bmpHeight;
  reg                 holdBuffer;
  wire                when_SuperResolutionPart1_l103;
  reg                 writeDone;
  wire                when_SuperResolutionPart1_l106;
  reg                 bufferRowCount_willIncrement;
  reg                 bufferRowCount_willClear;
  reg        [9:0]    bufferRowCount_valueNext;
  reg        [9:0]    bufferRowCount_value;
  wire                bufferRowCount_willOverflowIfInc;
  wire                bufferRowCount_willOverflow;
  reg                 bufferEnable;
  wire                when_SuperResolutionPart1_l112;
  wire                when_SuperResolutionPart1_l112_1;
  reg                 bufferSwitch;
  wire                when_SuperResolutionPart1_l115;
  reg                 nextRowBuffer;
  wire                when_SuperResolutionPart1_l118;
  reg                 bufferReuse;
  reg                 bufferWAddr_willIncrement;
  reg                 bufferWAddr_willClear;
  reg        [9:0]    bufferWAddr_valueNext;
  reg        [9:0]    bufferWAddr_value;
  wire                bufferWAddr_willOverflowIfInc;
  wire                bufferWAddr_willOverflow;
  reg                 outPixelAddr_willIncrement;
  reg                 outPixelAddr_willClear;
  reg        [10:0]   outPixelAddr_valueNext;
  reg        [10:0]   outPixelAddr_value;
  wire                outPixelAddr_willOverflowIfInc;
  wire                outPixelAddr_willOverflow;
  reg                 outRowCount_willIncrement;
  reg                 outRowCount_willClear;
  reg        [10:0]   outRowCount_valueNext;
  reg        [10:0]   outRowCount_value;
  wire                outRowCount_willOverflowIfInc;
  wire                outRowCount_willOverflow;
  reg                 outReachRowEnd;
  reg                 outReachFinalRow;
  reg                 bufferReachRowEnd;
  reg                 bufferReachFinalRow;
  reg        [9:0]    mainAddrOne;
  reg        [9:0]    counterAddrOne;
  reg        [9:0]    mainAddrTwo;
  reg        [9:0]    counterAddrTwo;
  wire                validStream_valid;
  reg                 validStream_ready;
  wire                controlStream_valid;
  wire                controlStream_ready;
  wire                controlStream_payload_frameStart;
  wire                controlStream_payload_rowEnd;
  wire                controlStream_payload_passMode;
  wire                controlStream_payload_passValid;
  wire       [2:0]    controlStream_payload_onceMode;
  wire                controlStream_payload_onceValid;
  wire                controlStream_payload_mainCompare;
  wire                controlStream_payload_counterCompare;
  wire       [7:0]    controlStream_payload_mainDiff;
  wire       [7:0]    controlStream_payload_counterDiff;
  wire                controlStream_payload_twiceCompValid;
  wire       [2:0]    controlStream_payload_twiceMode;
  reg                 controls_frameStart;
  reg                 controls_rowEnd;
  reg                 controls_passMode;
  reg                 controls_passValid;
  reg        [2:0]    controls_onceMode;
  reg                 controls_onceValid;
  wire                controls_mainCompare;
  wire                controls_counterCompare;
  wire       [7:0]    controls_mainDiff;
  wire       [7:0]    controls_counterDiff;
  reg                 controls_twiceCompValid;
  reg        [2:0]    controls_twiceMode;
  wire       [29:0]   CICC1851_controls_frameStart;
  wire                mainAddrOneStream_valid;
  wire                mainAddrOneStream_ready;
  wire       [9:0]    mainAddrOneStream_payload;
  wire                counterAddrOneStream_valid;
  wire                counterAddrOneStream_ready;
  wire       [9:0]    counterAddrOneStream_payload;
  wire                mainAddrTwoStream_valid;
  wire                mainAddrTwoStream_ready;
  wire       [9:0]    mainAddrTwoStream_payload;
  wire                counterAddrTwoStream_valid;
  wire                counterAddrTwoStream_ready;
  wire       [9:0]    counterAddrTwoStream_payload;
  wire                mainAddrOneStream_s2mPipe_valid;
  reg                 mainAddrOneStream_s2mPipe_ready;
  wire       [9:0]    mainAddrOneStream_s2mPipe_payload;
  reg                 mainAddrOneStream_rValid;
  reg        [9:0]    mainAddrOneStream_rData;
  wire                mainAddrOneStream_s2mPipe_m2sPipe_valid;
  wire                mainAddrOneStream_s2mPipe_m2sPipe_ready;
  wire       [9:0]    mainAddrOneStream_s2mPipe_m2sPipe_payload;
  reg                 mainAddrOneStream_s2mPipe_rValid;
  reg        [9:0]    mainAddrOneStream_s2mPipe_rData;
  wire                when_Stream_l368;
  wire                CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_mainOnePixelStream_payload;
  reg                 CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_1;
  reg                 CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_mainOnePixelStream_payload_1;
  wire                readStage_mainOnePixelStream_valid;
  wire                readStage_mainOnePixelStream_ready;
  wire       [7:0]    readStage_mainOnePixelStream_payload;
  reg                 CICC1851_readStage_mainOnePixelStream_valid;
  reg        [7:0]    CICC1851_readStage_mainOnePixelStream_payload_2;
  wire                when_Stream_l368_1;
  wire                counterAddrOneStream_s2mPipe_valid;
  reg                 counterAddrOneStream_s2mPipe_ready;
  wire       [9:0]    counterAddrOneStream_s2mPipe_payload;
  reg                 counterAddrOneStream_rValid;
  reg        [9:0]    counterAddrOneStream_rData;
  wire                counterAddrOneStream_s2mPipe_m2sPipe_valid;
  wire                counterAddrOneStream_s2mPipe_m2sPipe_ready;
  wire       [9:0]    counterAddrOneStream_s2mPipe_m2sPipe_payload;
  reg                 counterAddrOneStream_s2mPipe_rValid;
  reg        [9:0]    counterAddrOneStream_s2mPipe_rData;
  wire                when_Stream_l368_2;
  wire                CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_counterOnePixelStream_payload;
  reg                 CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_2;
  reg                 CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_counterOnePixelStream_payload_1;
  wire                readStage_counterOnePixelStream_valid;
  wire                readStage_counterOnePixelStream_ready;
  wire       [7:0]    readStage_counterOnePixelStream_payload;
  reg                 CICC1851_readStage_counterOnePixelStream_valid;
  reg        [7:0]    CICC1851_readStage_counterOnePixelStream_payload_2;
  wire                when_Stream_l368_3;
  wire                mainAddrTwoStream_s2mPipe_valid;
  reg                 mainAddrTwoStream_s2mPipe_ready;
  wire       [9:0]    mainAddrTwoStream_s2mPipe_payload;
  reg                 mainAddrTwoStream_rValid;
  reg        [9:0]    mainAddrTwoStream_rData;
  wire                mainAddrTwoStream_s2mPipe_m2sPipe_valid;
  wire                mainAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire       [9:0]    mainAddrTwoStream_s2mPipe_m2sPipe_payload;
  reg                 mainAddrTwoStream_s2mPipe_rValid;
  reg        [9:0]    mainAddrTwoStream_s2mPipe_rData;
  wire                when_Stream_l368_4;
  wire                CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_mainTwoPixelStream_payload;
  reg                 CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_3;
  reg                 CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_mainTwoPixelStream_payload_1;
  wire                readStage_mainTwoPixelStream_valid;
  wire                readStage_mainTwoPixelStream_ready;
  wire       [7:0]    readStage_mainTwoPixelStream_payload;
  reg                 CICC1851_readStage_mainTwoPixelStream_valid;
  reg        [7:0]    CICC1851_readStage_mainTwoPixelStream_payload_2;
  wire                when_Stream_l368_5;
  wire                counterAddrTwoStream_s2mPipe_valid;
  reg                 counterAddrTwoStream_s2mPipe_ready;
  wire       [9:0]    counterAddrTwoStream_s2mPipe_payload;
  reg                 counterAddrTwoStream_rValid;
  reg        [9:0]    counterAddrTwoStream_rData;
  wire                counterAddrTwoStream_s2mPipe_m2sPipe_valid;
  wire                counterAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire       [9:0]    counterAddrTwoStream_s2mPipe_m2sPipe_payload;
  reg                 counterAddrTwoStream_s2mPipe_rValid;
  reg        [9:0]    counterAddrTwoStream_s2mPipe_rData;
  wire                when_Stream_l368_6;
  wire                CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_counterTwoPixelStream_payload;
  reg                 CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_4;
  reg                 CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_counterTwoPixelStream_payload_1;
  wire                readStage_counterTwoPixelStream_valid;
  wire                readStage_counterTwoPixelStream_ready;
  wire       [7:0]    readStage_counterTwoPixelStream_payload;
  reg                 CICC1851_readStage_counterTwoPixelStream_valid;
  reg        [7:0]    CICC1851_readStage_counterTwoPixelStream_payload_2;
  wire                when_Stream_l368_7;
  wire                controlStream_s2mPipe_valid;
  reg                 controlStream_s2mPipe_ready;
  wire                controlStream_s2mPipe_payload_frameStart;
  wire                controlStream_s2mPipe_payload_rowEnd;
  wire                controlStream_s2mPipe_payload_passMode;
  wire                controlStream_s2mPipe_payload_passValid;
  wire       [2:0]    controlStream_s2mPipe_payload_onceMode;
  wire                controlStream_s2mPipe_payload_onceValid;
  wire                controlStream_s2mPipe_payload_mainCompare;
  wire                controlStream_s2mPipe_payload_counterCompare;
  wire       [7:0]    controlStream_s2mPipe_payload_mainDiff;
  wire       [7:0]    controlStream_s2mPipe_payload_counterDiff;
  wire                controlStream_s2mPipe_payload_twiceCompValid;
  wire       [2:0]    controlStream_s2mPipe_payload_twiceMode;
  reg                 controlStream_rValid;
  reg                 controlStream_rData_frameStart;
  reg                 controlStream_rData_rowEnd;
  reg                 controlStream_rData_passMode;
  reg                 controlStream_rData_passValid;
  reg        [2:0]    controlStream_rData_onceMode;
  reg                 controlStream_rData_onceValid;
  reg                 controlStream_rData_mainCompare;
  reg                 controlStream_rData_counterCompare;
  reg        [7:0]    controlStream_rData_mainDiff;
  reg        [7:0]    controlStream_rData_counterDiff;
  reg                 controlStream_rData_twiceCompValid;
  reg        [2:0]    controlStream_rData_twiceMode;
  wire                controlStream_s2mPipe_m2sPipe_valid;
  reg                 controlStream_s2mPipe_m2sPipe_ready;
  wire                controlStream_s2mPipe_m2sPipe_payload_frameStart;
  wire                controlStream_s2mPipe_m2sPipe_payload_rowEnd;
  wire                controlStream_s2mPipe_m2sPipe_payload_passMode;
  wire                controlStream_s2mPipe_m2sPipe_payload_passValid;
  wire       [2:0]    controlStream_s2mPipe_m2sPipe_payload_onceMode;
  wire                controlStream_s2mPipe_m2sPipe_payload_onceValid;
  wire                controlStream_s2mPipe_m2sPipe_payload_mainCompare;
  wire                controlStream_s2mPipe_m2sPipe_payload_counterCompare;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_payload_mainDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_payload_counterDiff;
  wire                controlStream_s2mPipe_m2sPipe_payload_twiceCompValid;
  wire       [2:0]    controlStream_s2mPipe_m2sPipe_payload_twiceMode;
  reg                 controlStream_s2mPipe_rValid;
  reg                 controlStream_s2mPipe_rData_frameStart;
  reg                 controlStream_s2mPipe_rData_rowEnd;
  reg                 controlStream_s2mPipe_rData_passMode;
  reg                 controlStream_s2mPipe_rData_passValid;
  reg        [2:0]    controlStream_s2mPipe_rData_onceMode;
  reg                 controlStream_s2mPipe_rData_onceValid;
  reg                 controlStream_s2mPipe_rData_mainCompare;
  reg                 controlStream_s2mPipe_rData_counterCompare;
  reg        [7:0]    controlStream_s2mPipe_rData_mainDiff;
  reg        [7:0]    controlStream_s2mPipe_rData_counterDiff;
  reg                 controlStream_s2mPipe_rData_twiceCompValid;
  reg        [2:0]    controlStream_s2mPipe_rData_twiceMode;
  wire                when_Stream_l368_8;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_valid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_ready;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_frameStart;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_rowEnd;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passMode;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passValid;
  wire       [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceMode;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceValid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainCompare;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterCompare;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDiff;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceCompValid;
  wire       [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceMode;
  reg                 controlStream_s2mPipe_m2sPipe_rValid;
  reg                 controlStream_s2mPipe_m2sPipe_rData_frameStart;
  reg                 controlStream_s2mPipe_m2sPipe_rData_rowEnd;
  reg                 controlStream_s2mPipe_m2sPipe_rData_passMode;
  reg                 controlStream_s2mPipe_m2sPipe_rData_passValid;
  reg        [2:0]    controlStream_s2mPipe_m2sPipe_rData_onceMode;
  reg                 controlStream_s2mPipe_m2sPipe_rData_onceValid;
  reg                 controlStream_s2mPipe_m2sPipe_rData_mainCompare;
  reg                 controlStream_s2mPipe_m2sPipe_rData_counterCompare;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_rData_mainDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_rData_counterDiff;
  reg                 controlStream_s2mPipe_m2sPipe_rData_twiceCompValid;
  reg        [2:0]    controlStream_s2mPipe_m2sPipe_rData_twiceMode;
  wire                when_Stream_l368_9;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_valid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_frameStart;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_rowEnd;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_passMode;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_passValid;
  wire       [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_onceMode;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_onceValid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainCompare;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterCompare;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterDiff;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_twiceCompValid;
  wire       [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_twiceMode;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_frameStart;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_rowEnd;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_passMode;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_passValid;
  reg        [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_onceMode;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_onceValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainCompare;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterCompare;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterDiff;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_twiceCompValid;
  reg        [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_twiceMode;
  wire                readStage_controlPipe_valid;
  wire                readStage_controlPipe_ready;
  wire                readStage_controlPipe_payload_frameStart;
  wire                readStage_controlPipe_payload_rowEnd;
  wire                readStage_controlPipe_payload_passMode;
  wire                readStage_controlPipe_payload_passValid;
  wire       [2:0]    readStage_controlPipe_payload_onceMode;
  wire                readStage_controlPipe_payload_onceValid;
  wire                readStage_controlPipe_payload_mainCompare;
  wire                readStage_controlPipe_payload_counterCompare;
  wire       [7:0]    readStage_controlPipe_payload_mainDiff;
  wire       [7:0]    readStage_controlPipe_payload_counterDiff;
  wire                readStage_controlPipe_payload_twiceCompValid;
  wire       [2:0]    readStage_controlPipe_payload_twiceMode;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_frameStart;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_rowEnd;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_passMode;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_passValid;
  reg        [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_onceMode;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_onceValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainCompare;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterCompare;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterDiff;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_twiceCompValid;
  reg        [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_twiceMode;
  wire                when_Stream_l368_10;
  wire                readStage_mainOnePixelStream_s2mPipe_valid;
  reg                 readStage_mainOnePixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_mainOnePixelStream_s2mPipe_payload;
  reg                 readStage_mainOnePixelStream_rValid;
  reg        [7:0]    readStage_mainOnePixelStream_rData;
  wire                compareStage_mainOnePixelStream_valid;
  wire                compareStage_mainOnePixelStream_ready;
  wire       [7:0]    compareStage_mainOnePixelStream_payload;
  reg                 readStage_mainOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_mainOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_11;
  wire                readStage_counterOnePixelStream_s2mPipe_valid;
  reg                 readStage_counterOnePixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_counterOnePixelStream_s2mPipe_payload;
  reg                 readStage_counterOnePixelStream_rValid;
  reg        [7:0]    readStage_counterOnePixelStream_rData;
  wire                compareStage_counterOnePixelStream_valid;
  wire                compareStage_counterOnePixelStream_ready;
  wire       [7:0]    compareStage_counterOnePixelStream_payload;
  reg                 readStage_counterOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_counterOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_12;
  wire                readStage_mainTwoPixelStream_s2mPipe_valid;
  reg                 readStage_mainTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_mainTwoPixelStream_s2mPipe_payload;
  reg                 readStage_mainTwoPixelStream_rValid;
  reg        [7:0]    readStage_mainTwoPixelStream_rData;
  wire                compareStage_mainTwoPixelStream_valid;
  wire                compareStage_mainTwoPixelStream_ready;
  wire       [7:0]    compareStage_mainTwoPixelStream_payload;
  reg                 readStage_mainTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_mainTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_13;
  wire                readStage_counterTwoPixelStream_s2mPipe_valid;
  reg                 readStage_counterTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_counterTwoPixelStream_s2mPipe_payload;
  reg                 readStage_counterTwoPixelStream_rValid;
  reg        [7:0]    readStage_counterTwoPixelStream_rData;
  wire                compareStage_counterTwoPixelStream_valid;
  wire                compareStage_counterTwoPixelStream_ready;
  wire       [7:0]    compareStage_counterTwoPixelStream_payload;
  reg                 readStage_counterTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_counterTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_14;
  reg                 CICC1851_readStage_controlPipe_translated_payload_mainCompare;
  reg                 CICC1851_readStage_controlPipe_translated_payload_counterCompare;
  wire                when_SuperResolutionPart1_l205;
  wire                when_SuperResolutionPart1_l209;
  wire                when_SuperResolutionPart1_l213;
  wire                when_SuperResolutionPart1_l217;
  wire                when_SuperResolutionPart1_l228;
  wire                when_SuperResolutionPart1_l230;
  wire                when_SuperResolutionPart1_l234;
  wire                when_SuperResolutionPart1_l236;
  wire                when_SuperResolutionPart1_l241;
  wire                when_SuperResolutionPart1_l246;
  wire                readStage_controlPipe_translated_valid;
  wire                readStage_controlPipe_translated_ready;
  wire                readStage_controlPipe_translated_payload_frameStart;
  wire                readStage_controlPipe_translated_payload_rowEnd;
  wire                readStage_controlPipe_translated_payload_passMode;
  wire                readStage_controlPipe_translated_payload_passValid;
  wire       [2:0]    readStage_controlPipe_translated_payload_onceMode;
  wire                readStage_controlPipe_translated_payload_onceValid;
  wire                readStage_controlPipe_translated_payload_mainCompare;
  wire                readStage_controlPipe_translated_payload_counterCompare;
  wire       [7:0]    readStage_controlPipe_translated_payload_mainDiff;
  wire       [7:0]    readStage_controlPipe_translated_payload_counterDiff;
  wire                readStage_controlPipe_translated_payload_twiceCompValid;
  wire       [2:0]    readStage_controlPipe_translated_payload_twiceMode;
  wire                readStage_controlPipe_translated_s2mPipe_valid;
  reg                 readStage_controlPipe_translated_s2mPipe_ready;
  wire                readStage_controlPipe_translated_s2mPipe_payload_frameStart;
  wire                readStage_controlPipe_translated_s2mPipe_payload_rowEnd;
  wire                readStage_controlPipe_translated_s2mPipe_payload_passMode;
  wire                readStage_controlPipe_translated_s2mPipe_payload_passValid;
  wire       [2:0]    readStage_controlPipe_translated_s2mPipe_payload_onceMode;
  wire                readStage_controlPipe_translated_s2mPipe_payload_onceValid;
  wire                readStage_controlPipe_translated_s2mPipe_payload_mainCompare;
  wire                readStage_controlPipe_translated_s2mPipe_payload_counterCompare;
  wire       [7:0]    readStage_controlPipe_translated_s2mPipe_payload_mainDiff;
  wire       [7:0]    readStage_controlPipe_translated_s2mPipe_payload_counterDiff;
  wire                readStage_controlPipe_translated_s2mPipe_payload_twiceCompValid;
  wire       [2:0]    readStage_controlPipe_translated_s2mPipe_payload_twiceMode;
  reg                 readStage_controlPipe_translated_rValid;
  reg                 readStage_controlPipe_translated_rData_frameStart;
  reg                 readStage_controlPipe_translated_rData_rowEnd;
  reg                 readStage_controlPipe_translated_rData_passMode;
  reg                 readStage_controlPipe_translated_rData_passValid;
  reg        [2:0]    readStage_controlPipe_translated_rData_onceMode;
  reg                 readStage_controlPipe_translated_rData_onceValid;
  reg                 readStage_controlPipe_translated_rData_mainCompare;
  reg                 readStage_controlPipe_translated_rData_counterCompare;
  reg        [7:0]    readStage_controlPipe_translated_rData_mainDiff;
  reg        [7:0]    readStage_controlPipe_translated_rData_counterDiff;
  reg                 readStage_controlPipe_translated_rData_twiceCompValid;
  reg        [2:0]    readStage_controlPipe_translated_rData_twiceMode;
  wire                compareStage_controlPipe_valid;
  wire                compareStage_controlPipe_ready;
  wire                compareStage_controlPipe_payload_frameStart;
  wire                compareStage_controlPipe_payload_rowEnd;
  wire                compareStage_controlPipe_payload_passMode;
  wire                compareStage_controlPipe_payload_passValid;
  wire       [2:0]    compareStage_controlPipe_payload_onceMode;
  wire                compareStage_controlPipe_payload_onceValid;
  wire                compareStage_controlPipe_payload_mainCompare;
  wire                compareStage_controlPipe_payload_counterCompare;
  wire       [7:0]    compareStage_controlPipe_payload_mainDiff;
  wire       [7:0]    compareStage_controlPipe_payload_counterDiff;
  wire                compareStage_controlPipe_payload_twiceCompValid;
  wire       [2:0]    compareStage_controlPipe_payload_twiceMode;
  reg                 readStage_controlPipe_translated_s2mPipe_rValid;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_frameStart;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_rowEnd;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_passMode;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_passValid;
  reg        [2:0]    readStage_controlPipe_translated_s2mPipe_rData_onceMode;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_onceValid;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_mainCompare;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_counterCompare;
  reg        [7:0]    readStage_controlPipe_translated_s2mPipe_rData_mainDiff;
  reg        [7:0]    readStage_controlPipe_translated_s2mPipe_rData_counterDiff;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_twiceCompValid;
  reg        [2:0]    readStage_controlPipe_translated_s2mPipe_rData_twiceMode;
  wire                when_Stream_l368_15;
  wire                compareStage_mainOnePixelStream_s2mPipe_valid;
  reg                 compareStage_mainOnePixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_mainOnePixelStream_s2mPipe_payload;
  reg                 compareStage_mainOnePixelStream_rValid;
  reg        [7:0]    compareStage_mainOnePixelStream_rData;
  wire                diffStage_mainOnePixelStream_valid;
  wire                diffStage_mainOnePixelStream_ready;
  wire       [7:0]    diffStage_mainOnePixelStream_payload;
  reg                 compareStage_mainOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_mainOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_16;
  wire                compareStage_counterOnePixelStream_s2mPipe_valid;
  reg                 compareStage_counterOnePixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_counterOnePixelStream_s2mPipe_payload;
  reg                 compareStage_counterOnePixelStream_rValid;
  reg        [7:0]    compareStage_counterOnePixelStream_rData;
  wire                diffStage_counterOnePixelStream_valid;
  wire                diffStage_counterOnePixelStream_ready;
  wire       [7:0]    diffStage_counterOnePixelStream_payload;
  reg                 compareStage_counterOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_counterOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_17;
  wire                compareStage_mainTwoPixelStream_s2mPipe_valid;
  reg                 compareStage_mainTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_mainTwoPixelStream_s2mPipe_payload;
  reg                 compareStage_mainTwoPixelStream_rValid;
  reg        [7:0]    compareStage_mainTwoPixelStream_rData;
  wire                diffStage_mainTwoPixelStream_valid;
  wire                diffStage_mainTwoPixelStream_ready;
  wire       [7:0]    diffStage_mainTwoPixelStream_payload;
  reg                 compareStage_mainTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_mainTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_18;
  wire                compareStage_counterTwoPixelStream_s2mPipe_valid;
  reg                 compareStage_counterTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_counterTwoPixelStream_s2mPipe_payload;
  reg                 compareStage_counterTwoPixelStream_rValid;
  reg        [7:0]    compareStage_counterTwoPixelStream_rData;
  wire                diffStage_counterTwoPixelStream_valid;
  wire                diffStage_counterTwoPixelStream_ready;
  wire       [7:0]    diffStage_counterTwoPixelStream_payload;
  reg                 compareStage_counterTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_counterTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_19;
  reg        [7:0]    CICC1851_compareStage_controlPipe_translated_payload_mainDiff;
  reg        [7:0]    CICC1851_compareStage_controlPipe_translated_payload_counterDiff;
  wire                compareStage_controlPipe_translated_valid;
  wire                compareStage_controlPipe_translated_ready;
  wire                compareStage_controlPipe_translated_payload_frameStart;
  wire                compareStage_controlPipe_translated_payload_rowEnd;
  wire                compareStage_controlPipe_translated_payload_passMode;
  wire                compareStage_controlPipe_translated_payload_passValid;
  wire       [2:0]    compareStage_controlPipe_translated_payload_onceMode;
  wire                compareStage_controlPipe_translated_payload_onceValid;
  wire                compareStage_controlPipe_translated_payload_mainCompare;
  wire                compareStage_controlPipe_translated_payload_counterCompare;
  wire       [7:0]    compareStage_controlPipe_translated_payload_mainDiff;
  wire       [7:0]    compareStage_controlPipe_translated_payload_counterDiff;
  wire                compareStage_controlPipe_translated_payload_twiceCompValid;
  wire       [2:0]    compareStage_controlPipe_translated_payload_twiceMode;
  wire                compareStage_controlPipe_translated_s2mPipe_valid;
  reg                 compareStage_controlPipe_translated_s2mPipe_ready;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_frameStart;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_rowEnd;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_passMode;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_passValid;
  wire       [2:0]    compareStage_controlPipe_translated_s2mPipe_payload_onceMode;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_onceValid;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_mainCompare;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_counterCompare;
  wire       [7:0]    compareStage_controlPipe_translated_s2mPipe_payload_mainDiff;
  wire       [7:0]    compareStage_controlPipe_translated_s2mPipe_payload_counterDiff;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_twiceCompValid;
  wire       [2:0]    compareStage_controlPipe_translated_s2mPipe_payload_twiceMode;
  reg                 compareStage_controlPipe_translated_rValid;
  reg                 compareStage_controlPipe_translated_rData_frameStart;
  reg                 compareStage_controlPipe_translated_rData_rowEnd;
  reg                 compareStage_controlPipe_translated_rData_passMode;
  reg                 compareStage_controlPipe_translated_rData_passValid;
  reg        [2:0]    compareStage_controlPipe_translated_rData_onceMode;
  reg                 compareStage_controlPipe_translated_rData_onceValid;
  reg                 compareStage_controlPipe_translated_rData_mainCompare;
  reg                 compareStage_controlPipe_translated_rData_counterCompare;
  reg        [7:0]    compareStage_controlPipe_translated_rData_mainDiff;
  reg        [7:0]    compareStage_controlPipe_translated_rData_counterDiff;
  reg                 compareStage_controlPipe_translated_rData_twiceCompValid;
  reg        [2:0]    compareStage_controlPipe_translated_rData_twiceMode;
  wire                diffStage_controlPipe_valid;
  wire                diffStage_controlPipe_ready;
  wire                diffStage_controlPipe_payload_frameStart;
  wire                diffStage_controlPipe_payload_rowEnd;
  wire                diffStage_controlPipe_payload_passMode;
  wire                diffStage_controlPipe_payload_passValid;
  wire       [2:0]    diffStage_controlPipe_payload_onceMode;
  wire                diffStage_controlPipe_payload_onceValid;
  wire                diffStage_controlPipe_payload_mainCompare;
  wire                diffStage_controlPipe_payload_counterCompare;
  wire       [7:0]    diffStage_controlPipe_payload_mainDiff;
  wire       [7:0]    diffStage_controlPipe_payload_counterDiff;
  wire                diffStage_controlPipe_payload_twiceCompValid;
  wire       [2:0]    diffStage_controlPipe_payload_twiceMode;
  reg                 compareStage_controlPipe_translated_s2mPipe_rValid;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_frameStart;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_rowEnd;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_passMode;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_passValid;
  reg        [2:0]    compareStage_controlPipe_translated_s2mPipe_rData_onceMode;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_onceValid;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_mainCompare;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_counterCompare;
  reg        [7:0]    compareStage_controlPipe_translated_s2mPipe_rData_mainDiff;
  reg        [7:0]    compareStage_controlPipe_translated_s2mPipe_rData_counterDiff;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_twiceCompValid;
  reg        [2:0]    compareStage_controlPipe_translated_s2mPipe_rData_twiceMode;
  wire                when_Stream_l368_20;
  wire                diffStage_mainOnePixelStream_s2mPipe_valid;
  reg                 diffStage_mainOnePixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_mainOnePixelStream_s2mPipe_payload;
  reg                 diffStage_mainOnePixelStream_rValid;
  reg        [7:0]    diffStage_mainOnePixelStream_rData;
  wire                resultStage_mainOnePixelStream_valid;
  wire                resultStage_mainOnePixelStream_ready;
  wire       [7:0]    resultStage_mainOnePixelStream_payload;
  reg                 diffStage_mainOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_mainOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_21;
  wire                diffStage_counterOnePixelStream_s2mPipe_valid;
  reg                 diffStage_counterOnePixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_counterOnePixelStream_s2mPipe_payload;
  reg                 diffStage_counterOnePixelStream_rValid;
  reg        [7:0]    diffStage_counterOnePixelStream_rData;
  wire                resultStage_counterOnePixelStream_valid;
  wire                resultStage_counterOnePixelStream_ready;
  wire       [7:0]    resultStage_counterOnePixelStream_payload;
  reg                 diffStage_counterOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_counterOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_22;
  wire                diffStage_mainTwoPixelStream_s2mPipe_valid;
  reg                 diffStage_mainTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_mainTwoPixelStream_s2mPipe_payload;
  reg                 diffStage_mainTwoPixelStream_rValid;
  reg        [7:0]    diffStage_mainTwoPixelStream_rData;
  wire                resultStage_mainTwoPixelStream_valid;
  wire                resultStage_mainTwoPixelStream_ready;
  wire       [7:0]    resultStage_mainTwoPixelStream_payload;
  reg                 diffStage_mainTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_mainTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_23;
  wire                diffStage_counterTwoPixelStream_s2mPipe_valid;
  reg                 diffStage_counterTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_counterTwoPixelStream_s2mPipe_payload;
  reg                 diffStage_counterTwoPixelStream_rValid;
  reg        [7:0]    diffStage_counterTwoPixelStream_rData;
  wire                resultStage_counterTwoPixelStream_valid;
  wire                resultStage_counterTwoPixelStream_ready;
  wire       [7:0]    resultStage_counterTwoPixelStream_payload;
  reg                 diffStage_counterTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_counterTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_24;
  wire                diffStage_controlPipe_fork_io_outputs_0_s2mPipe_valid;
  reg                 diffStage_controlPipe_fork_io_outputs_0_s2mPipe_ready;
  wire                diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_frameStart;
  wire                diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_rowEnd;
  wire                diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_passMode;
  wire                diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_passValid;
  wire       [2:0]    diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_onceMode;
  wire                diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_onceValid;
  wire                diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_mainCompare;
  wire                diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_counterCompare;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_mainDiff;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_counterDiff;
  wire                diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_twiceCompValid;
  wire       [2:0]    diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_twiceMode;
  reg                 diffStage_controlPipe_fork_io_outputs_0_rValid;
  reg                 diffStage_controlPipe_fork_io_outputs_0_rData_frameStart;
  reg                 diffStage_controlPipe_fork_io_outputs_0_rData_rowEnd;
  reg                 diffStage_controlPipe_fork_io_outputs_0_rData_passMode;
  reg                 diffStage_controlPipe_fork_io_outputs_0_rData_passValid;
  reg        [2:0]    diffStage_controlPipe_fork_io_outputs_0_rData_onceMode;
  reg                 diffStage_controlPipe_fork_io_outputs_0_rData_onceValid;
  reg                 diffStage_controlPipe_fork_io_outputs_0_rData_mainCompare;
  reg                 diffStage_controlPipe_fork_io_outputs_0_rData_counterCompare;
  reg        [7:0]    diffStage_controlPipe_fork_io_outputs_0_rData_mainDiff;
  reg        [7:0]    diffStage_controlPipe_fork_io_outputs_0_rData_counterDiff;
  reg                 diffStage_controlPipe_fork_io_outputs_0_rData_twiceCompValid;
  reg        [2:0]    diffStage_controlPipe_fork_io_outputs_0_rData_twiceMode;
  wire                resultStage_controlPipe_valid;
  wire                resultStage_controlPipe_ready;
  wire                resultStage_controlPipe_payload_frameStart;
  wire                resultStage_controlPipe_payload_rowEnd;
  wire                resultStage_controlPipe_payload_passMode;
  wire                resultStage_controlPipe_payload_passValid;
  wire       [2:0]    resultStage_controlPipe_payload_onceMode;
  wire                resultStage_controlPipe_payload_onceValid;
  wire                resultStage_controlPipe_payload_mainCompare;
  wire                resultStage_controlPipe_payload_counterCompare;
  wire       [7:0]    resultStage_controlPipe_payload_mainDiff;
  wire       [7:0]    resultStage_controlPipe_payload_counterDiff;
  wire                resultStage_controlPipe_payload_twiceCompValid;
  wire       [2:0]    resultStage_controlPipe_payload_twiceMode;
  reg                 diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rValid;
  reg                 diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_frameStart;
  reg                 diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_rowEnd;
  reg                 diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_passMode;
  reg                 diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_passValid;
  reg        [2:0]    diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_onceMode;
  reg                 diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_onceValid;
  reg                 diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_mainCompare;
  reg                 diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_counterCompare;
  reg        [7:0]    diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_mainDiff;
  reg        [7:0]    diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_counterDiff;
  reg                 diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_twiceCompValid;
  reg        [2:0]    diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_twiceMode;
  wire                when_Stream_l368_25;
  wire                resultStage_pixelStream_valid;
  wire                resultStage_pixelStream_ready;
  reg        [7:0]    resultStage_pixelStream_payload;
  wire                when_SuperResolutionPart1_l339;
  wire                when_SuperResolutionPart1_l343;
  wire                when_SuperResolutionPart1_l347;
  wire                when_SuperResolutionPart1_l351;
  wire                when_SuperResolutionPart1_l362;
  wire                when_SuperResolutionPart1_l363;
  wire                when_SuperResolutionPart1_l366;
  wire                when_SuperResolutionPart1_l371;
  wire                when_SuperResolutionPart1_l372;
  wire                when_SuperResolutionPart1_l375;
  wire                when_SuperResolutionPart1_l381;
  wire                when_SuperResolutionPart1_l386;
  wire                resultStage_pixelStream_s2mPipe_valid;
  reg                 resultStage_pixelStream_s2mPipe_ready;
  wire       [7:0]    resultStage_pixelStream_s2mPipe_payload;
  reg                 resultStage_pixelStream_rValid;
  reg        [7:0]    resultStage_pixelStream_rData;
  wire                resultStage_resultStream_valid;
  wire                resultStage_resultStream_ready;
  wire       [7:0]    resultStage_resultStream_payload;
  reg                 resultStage_pixelStream_s2mPipe_rValid;
  reg        [7:0]    resultStage_pixelStream_s2mPipe_rData;
  wire                when_Stream_l368_26;
  wire                CICC1851_resultStage_mainOnePixelStream_ready;
  reg                 CICC1851_resultStage_mainOnePixelStream_ready_1;
  wire                CICC1851_resultStage_mainOnePixelStream_ready_2;
  wire                when_Stream_l438;
  reg                 resultsJoin_valid;
  wire                resultsJoin_ready;
  wire                pixelsStream_valid;
  wire                pixelsStream_ready;
  wire       [7:0]    pixelsStream_payload_pixel;
  wire                pixelsStream_payload_frameStart;
  wire                pixelsStream_payload_rowEnd;
  wire                pixelsStream_s2mPipe_valid;
  reg                 pixelsStream_s2mPipe_ready;
  wire       [7:0]    pixelsStream_s2mPipe_payload_pixel;
  wire                pixelsStream_s2mPipe_payload_frameStart;
  wire                pixelsStream_s2mPipe_payload_rowEnd;
  reg                 pixelsStream_rValid;
  reg        [7:0]    pixelsStream_rData_pixel;
  reg                 pixelsStream_rData_frameStart;
  reg                 pixelsStream_rData_rowEnd;
  wire                pixelsStream_s2mPipe_m2sPipe_valid;
  wire                pixelsStream_s2mPipe_m2sPipe_ready;
  wire       [7:0]    pixelsStream_s2mPipe_m2sPipe_payload_pixel;
  wire                pixelsStream_s2mPipe_m2sPipe_payload_frameStart;
  wire                pixelsStream_s2mPipe_m2sPipe_payload_rowEnd;
  reg                 pixelsStream_s2mPipe_rValid;
  reg        [7:0]    pixelsStream_s2mPipe_rData_pixel;
  reg                 pixelsStream_s2mPipe_rData_frameStart;
  reg                 pixelsStream_s2mPipe_rData_rowEnd;
  wire                when_Stream_l368_27;
  wire                pixelsIn_s2mPipe_valid;
  reg                 pixelsIn_s2mPipe_ready;
  wire       [7:0]    pixelsIn_s2mPipe_payload_pixel;
  wire                pixelsIn_s2mPipe_payload_frameStart;
  wire                pixelsIn_s2mPipe_payload_rowEnd;
  reg                 pixelsIn_rValid;
  reg        [7:0]    pixelsIn_rData_pixel;
  reg                 pixelsIn_rData_frameStart;
  reg                 pixelsIn_rData_rowEnd;
  wire                pixelsIn_s2mPipe_m2sPipe_valid;
  wire                pixelsIn_s2mPipe_m2sPipe_ready;
  wire       [7:0]    pixelsIn_s2mPipe_m2sPipe_payload_pixel;
  wire                pixelsIn_s2mPipe_m2sPipe_payload_frameStart;
  wire                pixelsIn_s2mPipe_m2sPipe_payload_rowEnd;
  reg                 pixelsIn_s2mPipe_rValid;
  reg        [7:0]    pixelsIn_s2mPipe_rData_pixel;
  reg                 pixelsIn_s2mPipe_rData_frameStart;
  reg                 pixelsIn_s2mPipe_rData_rowEnd;
  wire                when_Stream_l368_28;
  wire                passPixels_valid;
  wire                passPixels_ready;
  wire       [7:0]    passPixels_payload_pixel;
  wire                passPixels_payload_frameStart;
  wire                passPixels_payload_rowEnd;
  wire                passPixels_fire;
  wire                when_SuperResolutionPart1_l421;
  wire                passPixels_fire_1;
  wire                when_SuperResolutionPart1_l422;
  wire                passPixels_fire_2;
  wire                when_SuperResolutionPart1_l425;
  wire                passPixels_fire_3;
  wire                when_SuperResolutionPart1_l438;
  wire                passPixels_fire_4;
  wire                when_SuperResolutionPart1_l439;
  wire                when_SuperResolutionPart1_l442;
  wire                controlStream_fire;
  wire                when_SuperResolutionPart1_l447;
  wire                when_SuperResolutionPart1_l449;
  wire                passPixels_fire_5;
  wire                when_SuperResolutionPart1_l453;
  wire                passPixels_fire_6;
  wire                passPixels_fire_7;
  wire                passPixels_fire_8;
  wire                controlStateMachine_wantExit;
  reg                 controlStateMachine_wantStart;
  wire                controlStateMachine_wantKill;
  reg        [2:0]    controlStateMachine_stateReg;
  reg        [2:0]    controlStateMachine_stateNext;
  wire                when_SuperResolutionPart1_l482;
  wire                passPixels_fire_9;
  wire                when_SuperResolutionPart1_l484;
  wire                passPixels_fire_10;
  wire                when_SuperResolutionPart1_l489;
  wire                controlStream_fire_1;
  wire                when_SuperResolutionPart1_l498;
  wire                passPixels_fire_11;
  wire                when_SuperResolutionPart1_l500;
  wire                controlStream_fire_2;
  wire                when_SuperResolutionPart1_l507;
  wire                controlStream_fire_3;
  wire                when_SuperResolutionPart1_l510;
  wire                controlStream_fire_4;
  wire                when_SuperResolutionPart1_l511;
  wire                controlStream_fire_5;
  wire                when_SuperResolutionPart1_l513;
  wire                controlStream_fire_6;
  wire                when_SuperResolutionPart1_l537;
  wire                controlStream_fire_7;
  wire                when_SuperResolutionPart1_l542;
  wire                controlStream_fire_8;
  wire                passPixels_fire_12;
  wire                when_SuperResolutionPart1_l563;
  wire                controlStream_fire_9;
  wire                when_SuperResolutionPart1_l578;
  wire                controlStream_fire_10;
  wire                when_SuperResolutionPart1_l579;
  wire                controlStream_fire_11;
  wire                when_SuperResolutionPart1_l581;
  wire                controlStream_fire_12;
  wire                controlStream_fire_13;
  wire                when_SuperResolutionPart1_l612;
  wire                controlStream_fire_14;
  wire                when_SuperResolutionPart1_l664;
  wire                controlStream_fire_15;
  wire                when_SuperResolutionPart1_l665;
  wire                controlStream_fire_16;
  wire                when_SuperResolutionPart1_l667;
  wire                controlStream_fire_17;
  `ifndef SYNTHESIS
  reg [39:0] controlStateMachine_stateReg_string;
  reg [39:0] controlStateMachine_stateNext_string;
  `endif

  reg [7:0] lineBufferOne [0:959];
  reg [7:0] lineBufferTwo [0:959];

  assign CICC1851_bufferRowCount_valueNext_1 = bufferRowCount_willIncrement;
  assign CICC1851_bufferRowCount_valueNext = {9'd0, CICC1851_bufferRowCount_valueNext_1};
  assign CICC1851_bufferWAddr_valueNext_1 = bufferWAddr_willIncrement;
  assign CICC1851_bufferWAddr_valueNext = {9'd0, CICC1851_bufferWAddr_valueNext_1};
  assign CICC1851_outPixelAddr_valueNext_1 = outPixelAddr_willIncrement;
  assign CICC1851_outPixelAddr_valueNext = {10'd0, CICC1851_outPixelAddr_valueNext_1};
  assign CICC1851_outRowCount_valueNext_1 = outRowCount_willIncrement;
  assign CICC1851_outRowCount_valueNext = {10'd0, CICC1851_outRowCount_valueNext_1};
  assign CICC1851_mainAddrOne = (outPixelAddr_value / 2'b10);
  assign CICC1851_counterAddrOne = (outPixelAddr_value / 2'b10);
  assign CICC1851_mainAddrTwo = (outPixelAddr_value / 2'b10);
  assign CICC1851_counterAddrTwo = (outPixelAddr_value / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload = (CICC1851_resultStage_pixelStream_payload_1 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_1 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_2 = (CICC1851_resultStage_pixelStream_payload_3 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_3 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_4 = (CICC1851_resultStage_pixelStream_payload_5 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_5 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_mainTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_6 = (CICC1851_resultStage_pixelStream_payload_7 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_7 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_mainOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_8 = (CICC1851_resultStage_pixelStream_payload_9 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_9 = ({1'b0,diffStage_counterOnePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_10 = (CICC1851_resultStage_pixelStream_payload_11 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_11 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_mainTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_12 = (CICC1851_resultStage_pixelStream_payload_13 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_13 = ({1'b0,diffStage_counterOnePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_14 = (CICC1851_resultStage_pixelStream_payload_15 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_15 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_mainTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_16 = (CICC1851_resultStage_pixelStream_payload_17 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_17 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_18 = (CICC1851_resultStage_pixelStream_payload_19 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_19 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_when_SuperResolutionPart1_l421 = (bmpWidth - 10'h002);
  assign CICC1851_when_SuperResolutionPart1_l422 = (bmpHeight - 10'h002);
  assign CICC1851_when_SuperResolutionPart1_l447 = (outRowCount_value % 2'b10);
  assign CICC1851_when_SuperResolutionPart1_l482 = (outRowCount_value % 2'b10);
  assign CICC1851_when_SuperResolutionPart1_l484 = (outPixelAddr_value % 2'b10);
  assign CICC1851_when_SuperResolutionPart1_l489 = (outPixelAddr_value % 2'b10);
  assign CICC1851_when_SuperResolutionPart1_l498 = {1'd0, outRowCount_value};
  assign CICC1851_when_SuperResolutionPart1_l498_1 = (2'b10 * bufferRowCount_value);
  assign CICC1851_when_SuperResolutionPart1_l500 = (2'b10 * bufferWAddr_value);
  assign CICC1851_when_SuperResolutionPart1_l500_1 = ({1'b0,outPixelAddr_value} + CICC1851_when_SuperResolutionPart1_l500_2);
  assign CICC1851_when_SuperResolutionPart1_l500_3 = {1'b0,2'b10};
  assign CICC1851_when_SuperResolutionPart1_l500_2 = {9'd0, CICC1851_when_SuperResolutionPart1_l500_3};
  assign CICC1851_when_SuperResolutionPart1_l510 = {1'd0, outPixelAddr_value};
  assign CICC1851_when_SuperResolutionPart1_l510_1 = (CICC1851_when_SuperResolutionPart1_l510_2 - 12'h002);
  assign CICC1851_when_SuperResolutionPart1_l510_2 = (2'b10 * bmpWidth);
  assign CICC1851_when_SuperResolutionPart1_l511 = {1'd0, outRowCount_value};
  assign CICC1851_when_SuperResolutionPart1_l511_1 = (CICC1851_when_SuperResolutionPart1_l511_2 - 12'h002);
  assign CICC1851_when_SuperResolutionPart1_l511_2 = (2'b10 * bmpHeight);
  assign CICC1851_when_SuperResolutionPart1_l537 = (outRowCount_value % 2'b10);
  assign CICC1851_when_SuperResolutionPart1_l542_1 = (11'h002 + outRowCount_value);
  assign CICC1851_when_SuperResolutionPart1_l542 = {1'd0, CICC1851_when_SuperResolutionPart1_l542_1};
  assign CICC1851_when_SuperResolutionPart1_l542_2 = (2'b10 * bufferRowCount_value);
  assign CICC1851_mainAddrOne_1 = (CICC1851_mainAddrOne_2 / 2'b10);
  assign CICC1851_mainAddrOne_2 = (outPixelAddr_value - 11'h001);
  assign CICC1851_counterAddrOne_1 = (CICC1851_counterAddrOne_2 / 2'b10);
  assign CICC1851_counterAddrOne_2 = (outPixelAddr_value - 11'h001);
  assign CICC1851_counterAddrOne_3 = (CICC1851_counterAddrOne_4 / 2'b10);
  assign CICC1851_counterAddrOne_4 = ({1'b0,outPixelAddr_value} + CICC1851_counterAddrOne_5);
  assign CICC1851_counterAddrOne_6 = {1'b0,1'b1};
  assign CICC1851_counterAddrOne_5 = {10'd0, CICC1851_counterAddrOne_6};
  assign CICC1851_controls_onceMode = 1'b1;
  assign CICC1851_mainAddrTwo_1 = (CICC1851_mainAddrTwo_2 / 2'b10);
  assign CICC1851_mainAddrTwo_2 = (outPixelAddr_value - 11'h001);
  assign CICC1851_counterAddrTwo_1 = (CICC1851_counterAddrTwo_2 / 2'b10);
  assign CICC1851_counterAddrTwo_2 = (outPixelAddr_value - 11'h001);
  assign CICC1851_counterAddrTwo_3 = (CICC1851_counterAddrTwo_4 / 2'b10);
  assign CICC1851_counterAddrTwo_4 = ({1'b0,outPixelAddr_value} + CICC1851_counterAddrTwo_5);
  assign CICC1851_counterAddrTwo_6 = {1'b0,1'b1};
  assign CICC1851_counterAddrTwo_5 = {10'd0, CICC1851_counterAddrTwo_6};
  assign CICC1851_when_SuperResolutionPart1_l563 = (2'b10 * bufferWAddr_value);
  assign CICC1851_when_SuperResolutionPart1_l563_1 = ({1'b0,outPixelAddr_value} + CICC1851_when_SuperResolutionPart1_l563_2);
  assign CICC1851_when_SuperResolutionPart1_l563_3 = {1'b0,2'b10};
  assign CICC1851_when_SuperResolutionPart1_l563_2 = {9'd0, CICC1851_when_SuperResolutionPart1_l563_3};
  assign CICC1851_controls_onceMode_1 = 2'b10;
  assign CICC1851_controls_onceMode_2 = 2'b11;
  assign CICC1851_mainAddrOne_3 = (outPixelAddr_value / 2'b10);
  assign CICC1851_mainAddrTwo_3 = (outPixelAddr_value / 2'b10);
  assign CICC1851_when_SuperResolutionPart1_l578 = {1'd0, outPixelAddr_value};
  assign CICC1851_when_SuperResolutionPart1_l578_1 = (CICC1851_when_SuperResolutionPart1_l578_2 - 12'h002);
  assign CICC1851_when_SuperResolutionPart1_l578_2 = (2'b10 * bmpWidth);
  assign CICC1851_when_SuperResolutionPart1_l579 = {1'd0, outRowCount_value};
  assign CICC1851_when_SuperResolutionPart1_l579_1 = (CICC1851_when_SuperResolutionPart1_l579_2 - 12'h002);
  assign CICC1851_when_SuperResolutionPart1_l579_2 = (2'b10 * bmpHeight);
  assign CICC1851_mainAddrOne_4 = (CICC1851_mainAddrOne_5 / 2'b10);
  assign CICC1851_mainAddrOne_5 = (outPixelAddr_value - 11'h001);
  assign CICC1851_mainAddrOne_6 = (CICC1851_mainAddrOne_7 / 2'b10);
  assign CICC1851_mainAddrOne_7 = (outPixelAddr_value - 11'h001);
  assign CICC1851_counterAddrOne_7 = (CICC1851_counterAddrOne_8 / 2'b10);
  assign CICC1851_counterAddrOne_8 = ({1'b0,outPixelAddr_value} + CICC1851_counterAddrOne_9);
  assign CICC1851_counterAddrOne_10 = {1'b0,1'b1};
  assign CICC1851_counterAddrOne_9 = {10'd0, CICC1851_counterAddrOne_10};
  assign CICC1851_mainAddrTwo_4 = (CICC1851_mainAddrTwo_5 / 2'b10);
  assign CICC1851_mainAddrTwo_5 = (outPixelAddr_value - 11'h001);
  assign CICC1851_mainAddrTwo_6 = (CICC1851_mainAddrTwo_7 / 2'b10);
  assign CICC1851_mainAddrTwo_7 = (outPixelAddr_value - 11'h001);
  assign CICC1851_counterAddrTwo_7 = (CICC1851_counterAddrTwo_8 / 2'b10);
  assign CICC1851_counterAddrTwo_8 = ({1'b0,outPixelAddr_value} + CICC1851_counterAddrTwo_9);
  assign CICC1851_counterAddrTwo_10 = {1'b0,1'b1};
  assign CICC1851_counterAddrTwo_9 = {10'd0, CICC1851_counterAddrTwo_10};
  assign CICC1851_mainAddrOne_8 = (CICC1851_mainAddrOne_9 / 2'b10);
  assign CICC1851_mainAddrOne_9 = (outPixelAddr_value - 11'h001);
  assign CICC1851_counterAddrTwo_11 = (CICC1851_counterAddrTwo_12 / 2'b10);
  assign CICC1851_counterAddrTwo_12 = (outPixelAddr_value - 11'h001);
  assign CICC1851_mainAddrTwo_8 = (CICC1851_mainAddrTwo_9 / 2'b10);
  assign CICC1851_mainAddrTwo_9 = (outPixelAddr_value - 11'h001);
  assign CICC1851_counterAddrOne_11 = (CICC1851_counterAddrOne_12 / 2'b10);
  assign CICC1851_counterAddrOne_12 = (outPixelAddr_value - 11'h001);
  assign CICC1851_mainAddrTwo_10 = (CICC1851_mainAddrTwo_11 / 2'b10);
  assign CICC1851_mainAddrTwo_11 = ({1'b0,outPixelAddr_value} + CICC1851_mainAddrTwo_12);
  assign CICC1851_mainAddrTwo_13 = {1'b0,1'b1};
  assign CICC1851_mainAddrTwo_12 = {10'd0, CICC1851_mainAddrTwo_13};
  assign CICC1851_counterAddrOne_13 = (CICC1851_counterAddrOne_14 / 2'b10);
  assign CICC1851_counterAddrOne_14 = ({1'b0,outPixelAddr_value} + CICC1851_counterAddrOne_15);
  assign CICC1851_counterAddrOne_16 = {1'b0,1'b1};
  assign CICC1851_counterAddrOne_15 = {10'd0, CICC1851_counterAddrOne_16};
  assign CICC1851_mainAddrTwo_14 = (CICC1851_mainAddrTwo_15 / 2'b10);
  assign CICC1851_mainAddrTwo_15 = (outPixelAddr_value - 11'h001);
  assign CICC1851_counterAddrOne_17 = (CICC1851_counterAddrOne_18 / 2'b10);
  assign CICC1851_counterAddrOne_18 = (outPixelAddr_value - 11'h001);
  assign CICC1851_mainAddrOne_10 = (CICC1851_mainAddrOne_11 / 2'b10);
  assign CICC1851_mainAddrOne_11 = (outPixelAddr_value - 11'h001);
  assign CICC1851_counterAddrTwo_13 = (CICC1851_counterAddrTwo_14 / 2'b10);
  assign CICC1851_counterAddrTwo_14 = (outPixelAddr_value - 11'h001);
  assign CICC1851_mainAddrOne_12 = (CICC1851_mainAddrOne_13 / 2'b10);
  assign CICC1851_mainAddrOne_13 = ({1'b0,outPixelAddr_value} + CICC1851_mainAddrOne_14);
  assign CICC1851_mainAddrOne_15 = {1'b0,1'b1};
  assign CICC1851_mainAddrOne_14 = {10'd0, CICC1851_mainAddrOne_15};
  assign CICC1851_counterAddrTwo_15 = (CICC1851_counterAddrTwo_16 / 2'b10);
  assign CICC1851_counterAddrTwo_16 = ({1'b0,outPixelAddr_value} + CICC1851_counterAddrTwo_17);
  assign CICC1851_counterAddrTwo_18 = {1'b0,1'b1};
  assign CICC1851_counterAddrTwo_17 = {10'd0, CICC1851_counterAddrTwo_18};
  assign CICC1851_when_SuperResolutionPart1_l664 = {1'd0, outPixelAddr_value};
  assign CICC1851_when_SuperResolutionPart1_l664_1 = (CICC1851_when_SuperResolutionPart1_l664_2 - 12'h002);
  assign CICC1851_when_SuperResolutionPart1_l664_2 = (2'b10 * bmpWidth);
  assign CICC1851_when_SuperResolutionPart1_l665 = {1'd0, outRowCount_value};
  assign CICC1851_when_SuperResolutionPart1_l665_1 = (CICC1851_when_SuperResolutionPart1_l665_2 - 12'h002);
  assign CICC1851_when_SuperResolutionPart1_l665_2 = (2'b10 * bmpHeight);
  assign CICC1851_lineBufferOne_port = passPixels_payload_pixel;
  assign CICC1851_lineBufferOne_port_1 = (passPixels_fire_7 && (! bufferSwitch));
  assign CICC1851_lineBufferTwo_port = passPixels_payload_pixel;
  assign CICC1851_lineBufferTwo_port_1 = (passPixels_fire_6 && bufferSwitch);
  always @(posedge clk) begin
    if(mainAddrOneStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferOne_port0 <= lineBufferOne[mainAddrOneStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(counterAddrOneStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferOne_port1 <= lineBufferOne[counterAddrOneStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(CICC1851_lineBufferOne_port_1) begin
      lineBufferOne[bufferWAddr_value] <= CICC1851_lineBufferOne_port;
    end
  end

  always @(posedge clk) begin
    if(mainAddrTwoStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferTwo_port0 <= lineBufferTwo[mainAddrTwoStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(counterAddrTwoStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferTwo_port1 <= lineBufferTwo[counterAddrTwoStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(CICC1851_lineBufferTwo_port_1) begin
      lineBufferTwo[bufferWAddr_value] <= CICC1851_lineBufferTwo_port;
    end
  end

  StreamFork_1 diffStage_controlPipe_fork (
    .io_input_valid                      (diffStage_controlPipe_valid                                     ), //i
    .io_input_ready                      (diffStage_controlPipe_fork_io_input_ready                       ), //o
    .io_input_payload_frameStart         (diffStage_controlPipe_payload_frameStart                        ), //i
    .io_input_payload_rowEnd             (diffStage_controlPipe_payload_rowEnd                            ), //i
    .io_input_payload_passMode           (diffStage_controlPipe_payload_passMode                          ), //i
    .io_input_payload_passValid          (diffStage_controlPipe_payload_passValid                         ), //i
    .io_input_payload_onceMode           (diffStage_controlPipe_payload_onceMode[2:0]                     ), //i
    .io_input_payload_onceValid          (diffStage_controlPipe_payload_onceValid                         ), //i
    .io_input_payload_mainCompare        (diffStage_controlPipe_payload_mainCompare                       ), //i
    .io_input_payload_counterCompare     (diffStage_controlPipe_payload_counterCompare                    ), //i
    .io_input_payload_mainDiff           (diffStage_controlPipe_payload_mainDiff[7:0]                     ), //i
    .io_input_payload_counterDiff        (diffStage_controlPipe_payload_counterDiff[7:0]                  ), //i
    .io_input_payload_twiceCompValid     (diffStage_controlPipe_payload_twiceCompValid                    ), //i
    .io_input_payload_twiceMode          (diffStage_controlPipe_payload_twiceMode[2:0]                    ), //i
    .io_outputs_0_valid                  (diffStage_controlPipe_fork_io_outputs_0_valid                   ), //o
    .io_outputs_0_ready                  (diffStage_controlPipe_fork_io_outputs_0_ready                   ), //i
    .io_outputs_0_payload_frameStart     (diffStage_controlPipe_fork_io_outputs_0_payload_frameStart      ), //o
    .io_outputs_0_payload_rowEnd         (diffStage_controlPipe_fork_io_outputs_0_payload_rowEnd          ), //o
    .io_outputs_0_payload_passMode       (diffStage_controlPipe_fork_io_outputs_0_payload_passMode        ), //o
    .io_outputs_0_payload_passValid      (diffStage_controlPipe_fork_io_outputs_0_payload_passValid       ), //o
    .io_outputs_0_payload_onceMode       (diffStage_controlPipe_fork_io_outputs_0_payload_onceMode[2:0]   ), //o
    .io_outputs_0_payload_onceValid      (diffStage_controlPipe_fork_io_outputs_0_payload_onceValid       ), //o
    .io_outputs_0_payload_mainCompare    (diffStage_controlPipe_fork_io_outputs_0_payload_mainCompare     ), //o
    .io_outputs_0_payload_counterCompare (diffStage_controlPipe_fork_io_outputs_0_payload_counterCompare  ), //o
    .io_outputs_0_payload_mainDiff       (diffStage_controlPipe_fork_io_outputs_0_payload_mainDiff[7:0]   ), //o
    .io_outputs_0_payload_counterDiff    (diffStage_controlPipe_fork_io_outputs_0_payload_counterDiff[7:0]), //o
    .io_outputs_0_payload_twiceCompValid (diffStage_controlPipe_fork_io_outputs_0_payload_twiceCompValid  ), //o
    .io_outputs_0_payload_twiceMode      (diffStage_controlPipe_fork_io_outputs_0_payload_twiceMode[2:0]  ), //o
    .io_outputs_1_valid                  (diffStage_controlPipe_fork_io_outputs_1_valid                   ), //o
    .io_outputs_1_ready                  (resultStage_pixelStream_ready                                   ), //i
    .io_outputs_1_payload_frameStart     (diffStage_controlPipe_fork_io_outputs_1_payload_frameStart      ), //o
    .io_outputs_1_payload_rowEnd         (diffStage_controlPipe_fork_io_outputs_1_payload_rowEnd          ), //o
    .io_outputs_1_payload_passMode       (diffStage_controlPipe_fork_io_outputs_1_payload_passMode        ), //o
    .io_outputs_1_payload_passValid      (diffStage_controlPipe_fork_io_outputs_1_payload_passValid       ), //o
    .io_outputs_1_payload_onceMode       (diffStage_controlPipe_fork_io_outputs_1_payload_onceMode[2:0]   ), //o
    .io_outputs_1_payload_onceValid      (diffStage_controlPipe_fork_io_outputs_1_payload_onceValid       ), //o
    .io_outputs_1_payload_mainCompare    (diffStage_controlPipe_fork_io_outputs_1_payload_mainCompare     ), //o
    .io_outputs_1_payload_counterCompare (diffStage_controlPipe_fork_io_outputs_1_payload_counterCompare  ), //o
    .io_outputs_1_payload_mainDiff       (diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff[7:0]   ), //o
    .io_outputs_1_payload_counterDiff    (diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff[7:0]), //o
    .io_outputs_1_payload_twiceCompValid (diffStage_controlPipe_fork_io_outputs_1_payload_twiceCompValid  ), //o
    .io_outputs_1_payload_twiceMode      (diffStage_controlPipe_fork_io_outputs_1_payload_twiceMode[2:0]  )  //o
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_6_BOOT : controlStateMachine_stateReg_string = "BOOT ";
      controlStateMachine_enumDef_6_HOLD : controlStateMachine_stateReg_string = "HOLD ";
      controlStateMachine_enumDef_6_PASS : controlStateMachine_stateReg_string = "PASS ";
      controlStateMachine_enumDef_6_ONCE : controlStateMachine_stateReg_string = "ONCE ";
      controlStateMachine_enumDef_6_TWICE : controlStateMachine_stateReg_string = "TWICE";
      default : controlStateMachine_stateReg_string = "?????";
    endcase
  end
  always @(*) begin
    case(controlStateMachine_stateNext)
      controlStateMachine_enumDef_6_BOOT : controlStateMachine_stateNext_string = "BOOT ";
      controlStateMachine_enumDef_6_HOLD : controlStateMachine_stateNext_string = "HOLD ";
      controlStateMachine_enumDef_6_PASS : controlStateMachine_stateNext_string = "PASS ";
      controlStateMachine_enumDef_6_ONCE : controlStateMachine_stateNext_string = "ONCE ";
      controlStateMachine_enumDef_6_TWICE : controlStateMachine_stateNext_string = "TWICE";
      default : controlStateMachine_stateNext_string = "?????";
    endcase
  end
  `endif

  always @(*) begin
    pixelsIn_ready = 1'b0;
    pixelsIn_ready = (! pixelsIn_rValid);
  end

  always @(*) begin
    pixelsOut_valid = 1'b0;
    pixelsOut_valid = pixelsStream_s2mPipe_m2sPipe_valid;
  end

  always @(*) begin
    pixelsOut_payload_pixel = 8'h0;
    pixelsOut_payload_pixel = pixelsStream_s2mPipe_m2sPipe_payload_pixel;
  end

  always @(*) begin
    pixelsOut_payload_frameStart = 1'b0;
    pixelsOut_payload_frameStart = pixelsStream_s2mPipe_m2sPipe_payload_frameStart;
  end

  always @(*) begin
    pixelsOut_payload_rowEnd = 1'b0;
    pixelsOut_payload_rowEnd = pixelsStream_s2mPipe_m2sPipe_payload_rowEnd;
  end

  always @(*) begin
    startOut = 1'b0;
    startOut = slaveStart;
  end

  always @(*) begin
    inpDoneOut = 1'b0;
    inpDoneOut = inpDone;
  end

  assign when_SuperResolutionPart1_l79 = (inpThreeDoneIn && inpTwoDoneIn);
  assign when_SuperResolutionPart1_l79_1 = (startIn && (! startIn_regNext));
  assign when_SuperResolutionPart1_l82 = (! startIn);
  assign when_SuperResolutionPart1_l85 = (startIn && (! readDone));
  assign when_SuperResolutionPart1_l85_1 = (! startIn);
  assign pixelsIn_fire = (pixelsIn_valid && pixelsIn_ready);
  assign when_SuperResolutionPart1_l88 = ((! inpTwoDoneIn) && pixelsIn_fire);
  assign when_SuperResolutionPart1_l88_1 = ((inpTwoDoneIn && inpThreeDoneIn) || (! startIn));
  assign when_SuperResolutionPart1_l103 = (! startIn);
  assign when_SuperResolutionPart1_l106 = (! startIn);
  always @(*) begin
    bufferRowCount_willIncrement = 1'b0;
    if(when_SuperResolutionPart1_l425) begin
      if(!bufferReachFinalRow) begin
        bufferRowCount_willIncrement = 1'b1;
      end
    end
  end

  always @(*) begin
    bufferRowCount_willClear = 1'b0;
    if(when_SuperResolutionPart1_l425) begin
      if(bufferReachFinalRow) begin
        bufferRowCount_willClear = 1'b1;
      end
    end
  end

  assign bufferRowCount_willOverflowIfInc = (bufferRowCount_value == 10'h21c);
  assign bufferRowCount_willOverflow = (bufferRowCount_willOverflowIfInc && bufferRowCount_willIncrement);
  always @(*) begin
    if(bufferRowCount_willOverflow) begin
      bufferRowCount_valueNext = 10'h0;
    end else begin
      bufferRowCount_valueNext = (bufferRowCount_value + CICC1851_bufferRowCount_valueNext);
    end
    if(bufferRowCount_willClear) begin
      bufferRowCount_valueNext = 10'h0;
    end
  end

  assign when_SuperResolutionPart1_l112 = ((startIn && (! holdBuffer)) && (! writeDone));
  assign when_SuperResolutionPart1_l112_1 = (((! startIn) || holdBuffer) || writeDone);
  assign when_SuperResolutionPart1_l115 = (! startRead);
  assign when_SuperResolutionPart1_l118 = (! startRead);
  always @(*) begin
    bufferWAddr_willIncrement = 1'b0;
    if(passPixels_fire_8) begin
      if(!passPixels_payload_rowEnd) begin
        bufferWAddr_willIncrement = 1'b1;
      end
    end
  end

  always @(*) begin
    bufferWAddr_willClear = 1'b0;
    if(passPixels_fire_8) begin
      if(passPixels_payload_rowEnd) begin
        bufferWAddr_willClear = 1'b1;
      end
    end
  end

  assign bufferWAddr_willOverflowIfInc = (bufferWAddr_value == 10'h3bf);
  assign bufferWAddr_willOverflow = (bufferWAddr_willOverflowIfInc && bufferWAddr_willIncrement);
  always @(*) begin
    if(bufferWAddr_willOverflow) begin
      bufferWAddr_valueNext = 10'h0;
    end else begin
      bufferWAddr_valueNext = (bufferWAddr_value + CICC1851_bufferWAddr_valueNext);
    end
    if(bufferWAddr_willClear) begin
      bufferWAddr_valueNext = 10'h0;
    end
  end

  always @(*) begin
    outPixelAddr_willIncrement = 1'b0;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_6_HOLD : begin
      end
      controlStateMachine_enumDef_6_PASS : begin
        if(controlStream_fire_6) begin
          if(!outReachRowEnd) begin
            outPixelAddr_willIncrement = 1'b1;
          end
        end
      end
      controlStateMachine_enumDef_6_ONCE : begin
        if(controlStream_fire_12) begin
          if(!outReachRowEnd) begin
            outPixelAddr_willIncrement = 1'b1;
          end
        end
      end
      controlStateMachine_enumDef_6_TWICE : begin
        if(controlStream_fire_17) begin
          if(!outReachRowEnd) begin
            outPixelAddr_willIncrement = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outPixelAddr_willClear = 1'b0;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_6_HOLD : begin
      end
      controlStateMachine_enumDef_6_PASS : begin
        if(controlStream_fire_6) begin
          if(outReachRowEnd) begin
            outPixelAddr_willClear = 1'b1;
          end
        end
      end
      controlStateMachine_enumDef_6_ONCE : begin
        if(controlStream_fire_12) begin
          if(outReachRowEnd) begin
            outPixelAddr_willClear = 1'b1;
          end
        end
      end
      controlStateMachine_enumDef_6_TWICE : begin
        if(controlStream_fire_17) begin
          if(outReachRowEnd) begin
            outPixelAddr_willClear = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign outPixelAddr_willOverflowIfInc = (outPixelAddr_value == 11'h77f);
  assign outPixelAddr_willOverflow = (outPixelAddr_willOverflowIfInc && outPixelAddr_willIncrement);
  always @(*) begin
    if(outPixelAddr_willOverflow) begin
      outPixelAddr_valueNext = 11'h0;
    end else begin
      outPixelAddr_valueNext = (outPixelAddr_value + CICC1851_outPixelAddr_valueNext);
    end
    if(outPixelAddr_willClear) begin
      outPixelAddr_valueNext = 11'h0;
    end
  end

  always @(*) begin
    outRowCount_willIncrement = 1'b0;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_6_HOLD : begin
      end
      controlStateMachine_enumDef_6_PASS : begin
        if(when_SuperResolutionPart1_l513) begin
          if(!outReachFinalRow) begin
            outRowCount_willIncrement = 1'b1;
          end
        end
      end
      controlStateMachine_enumDef_6_ONCE : begin
        if(when_SuperResolutionPart1_l581) begin
          if(!outReachFinalRow) begin
            outRowCount_willIncrement = 1'b1;
          end
        end
      end
      controlStateMachine_enumDef_6_TWICE : begin
        if(when_SuperResolutionPart1_l667) begin
          if(!outReachFinalRow) begin
            outRowCount_willIncrement = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outRowCount_willClear = 1'b0;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_6_HOLD : begin
      end
      controlStateMachine_enumDef_6_PASS : begin
        if(when_SuperResolutionPart1_l513) begin
          if(outReachFinalRow) begin
            outRowCount_willClear = 1'b1;
          end
        end
      end
      controlStateMachine_enumDef_6_ONCE : begin
        if(when_SuperResolutionPart1_l581) begin
          if(outReachFinalRow) begin
            outRowCount_willClear = 1'b1;
          end
        end
      end
      controlStateMachine_enumDef_6_TWICE : begin
        if(when_SuperResolutionPart1_l667) begin
          if(outReachFinalRow) begin
            outRowCount_willClear = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign outRowCount_willOverflowIfInc = (outRowCount_value == 11'h438);
  assign outRowCount_willOverflow = (outRowCount_willOverflowIfInc && outRowCount_willIncrement);
  always @(*) begin
    if(outRowCount_willOverflow) begin
      outRowCount_valueNext = 11'h0;
    end else begin
      outRowCount_valueNext = (outRowCount_value + CICC1851_outRowCount_valueNext);
    end
    if(outRowCount_willClear) begin
      outRowCount_valueNext = 11'h0;
    end
  end

  always @(*) begin
    mainAddrOne = CICC1851_mainAddrOne[9:0];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_6_HOLD : begin
      end
      controlStateMachine_enumDef_6_PASS : begin
      end
      controlStateMachine_enumDef_6_ONCE : begin
        if(when_SuperResolutionPart1_l537) begin
          if(nextRowBuffer) begin
            mainAddrOne = CICC1851_mainAddrOne_1[9:0];
          end
        end else begin
          mainAddrOne = CICC1851_mainAddrOne_3[9:0];
        end
      end
      controlStateMachine_enumDef_6_TWICE : begin
        if(outReachFinalRow) begin
          if(nextRowBuffer) begin
            if(outReachRowEnd) begin
              mainAddrOne = CICC1851_mainAddrOne_4[9:0];
            end else begin
              mainAddrOne = CICC1851_mainAddrOne_6[9:0];
            end
          end
        end else begin
          if(nextRowBuffer) begin
            mainAddrOne = CICC1851_mainAddrOne_8[9:0];
          end else begin
            if(outReachRowEnd) begin
              mainAddrOne = CICC1851_mainAddrOne_10[9:0];
            end else begin
              mainAddrOne = CICC1851_mainAddrOne_12[9:0];
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    counterAddrOne = CICC1851_counterAddrOne[9:0];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_6_HOLD : begin
      end
      controlStateMachine_enumDef_6_PASS : begin
      end
      controlStateMachine_enumDef_6_ONCE : begin
        if(when_SuperResolutionPart1_l537) begin
          if(nextRowBuffer) begin
            if(outReachRowEnd) begin
              counterAddrOne = CICC1851_counterAddrOne_1[9:0];
            end else begin
              counterAddrOne = CICC1851_counterAddrOne_3[9:0];
            end
          end
        end
      end
      controlStateMachine_enumDef_6_TWICE : begin
        if(outReachFinalRow) begin
          if(nextRowBuffer) begin
            if(!outReachRowEnd) begin
              counterAddrOne = CICC1851_counterAddrOne_7[9:0];
            end
          end
        end else begin
          if(nextRowBuffer) begin
            if(outReachRowEnd) begin
              counterAddrOne = CICC1851_counterAddrOne_11[9:0];
            end else begin
              counterAddrOne = CICC1851_counterAddrOne_13[9:0];
            end
          end else begin
            counterAddrOne = CICC1851_counterAddrOne_17[9:0];
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    mainAddrTwo = CICC1851_mainAddrTwo[9:0];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_6_HOLD : begin
      end
      controlStateMachine_enumDef_6_PASS : begin
      end
      controlStateMachine_enumDef_6_ONCE : begin
        if(when_SuperResolutionPart1_l537) begin
          if(!nextRowBuffer) begin
            mainAddrTwo = CICC1851_mainAddrTwo_1[9:0];
          end
        end else begin
          mainAddrTwo = CICC1851_mainAddrTwo_3[9:0];
        end
      end
      controlStateMachine_enumDef_6_TWICE : begin
        if(outReachFinalRow) begin
          if(!nextRowBuffer) begin
            if(outReachRowEnd) begin
              mainAddrTwo = CICC1851_mainAddrTwo_4[9:0];
            end else begin
              mainAddrTwo = CICC1851_mainAddrTwo_6[9:0];
            end
          end
        end else begin
          if(nextRowBuffer) begin
            if(outReachRowEnd) begin
              mainAddrTwo = CICC1851_mainAddrTwo_8[9:0];
            end else begin
              mainAddrTwo = CICC1851_mainAddrTwo_10[9:0];
            end
          end else begin
            mainAddrTwo = CICC1851_mainAddrTwo_14[9:0];
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    counterAddrTwo = CICC1851_counterAddrTwo[9:0];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_6_HOLD : begin
      end
      controlStateMachine_enumDef_6_PASS : begin
      end
      controlStateMachine_enumDef_6_ONCE : begin
        if(when_SuperResolutionPart1_l537) begin
          if(!nextRowBuffer) begin
            if(outReachRowEnd) begin
              counterAddrTwo = CICC1851_counterAddrTwo_1[9:0];
            end else begin
              counterAddrTwo = CICC1851_counterAddrTwo_3[9:0];
            end
          end
        end
      end
      controlStateMachine_enumDef_6_TWICE : begin
        if(outReachFinalRow) begin
          if(!nextRowBuffer) begin
            if(!outReachRowEnd) begin
              counterAddrTwo = CICC1851_counterAddrTwo_7[9:0];
            end
          end
        end else begin
          if(nextRowBuffer) begin
            counterAddrTwo = CICC1851_counterAddrTwo_11[9:0];
          end else begin
            if(outReachRowEnd) begin
              counterAddrTwo = CICC1851_counterAddrTwo_13[9:0];
            end else begin
              counterAddrTwo = CICC1851_counterAddrTwo_15[9:0];
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign validStream_valid = 1'b1;
  assign CICC1851_controls_frameStart = 30'h0;
  always @(*) begin
    controls_frameStart = CICC1851_controls_frameStart[0];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_6_HOLD : begin
      end
      controlStateMachine_enumDef_6_PASS : begin
        if(frameStart) begin
          controls_frameStart = 1'b1;
        end
      end
      controlStateMachine_enumDef_6_ONCE : begin
      end
      controlStateMachine_enumDef_6_TWICE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_rowEnd = CICC1851_controls_frameStart[1];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_6_HOLD : begin
      end
      controlStateMachine_enumDef_6_PASS : begin
        if(outReachRowEnd) begin
          controls_rowEnd = 1'b1;
        end
      end
      controlStateMachine_enumDef_6_ONCE : begin
        if(outReachRowEnd) begin
          controls_rowEnd = 1'b1;
        end
      end
      controlStateMachine_enumDef_6_TWICE : begin
        if(outReachRowEnd) begin
          controls_rowEnd = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_passMode = CICC1851_controls_frameStart[2];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_6_HOLD : begin
      end
      controlStateMachine_enumDef_6_PASS : begin
        if(nextRowBuffer) begin
          controls_passMode = 1'b0;
        end else begin
          controls_passMode = 1'b1;
        end
      end
      controlStateMachine_enumDef_6_ONCE : begin
      end
      controlStateMachine_enumDef_6_TWICE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_passValid = CICC1851_controls_frameStart[3];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_6_HOLD : begin
      end
      controlStateMachine_enumDef_6_PASS : begin
        controls_passValid = 1'b1;
      end
      controlStateMachine_enumDef_6_ONCE : begin
      end
      controlStateMachine_enumDef_6_TWICE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_onceMode = CICC1851_controls_frameStart[6 : 4];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_6_HOLD : begin
      end
      controlStateMachine_enumDef_6_PASS : begin
      end
      controlStateMachine_enumDef_6_ONCE : begin
        if(when_SuperResolutionPart1_l537) begin
          if(nextRowBuffer) begin
            controls_onceMode = 3'b000;
          end else begin
            controls_onceMode = {2'd0, CICC1851_controls_onceMode};
          end
        end else begin
          if(outReachFinalRow) begin
            if(nextRowBuffer) begin
              controls_onceMode = 3'b101;
            end else begin
              controls_onceMode = 3'b100;
            end
          end else begin
            if(nextRowBuffer) begin
              controls_onceMode = {1'd0, CICC1851_controls_onceMode_1};
            end else begin
              controls_onceMode = {1'd0, CICC1851_controls_onceMode_2};
            end
          end
        end
      end
      controlStateMachine_enumDef_6_TWICE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_onceValid = CICC1851_controls_frameStart[7];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_6_HOLD : begin
      end
      controlStateMachine_enumDef_6_PASS : begin
      end
      controlStateMachine_enumDef_6_ONCE : begin
        controls_onceValid = 1'b1;
      end
      controlStateMachine_enumDef_6_TWICE : begin
      end
      default : begin
      end
    endcase
  end

  assign controls_mainCompare = CICC1851_controls_frameStart[8];
  assign controls_counterCompare = CICC1851_controls_frameStart[9];
  assign controls_mainDiff = CICC1851_controls_frameStart[17 : 10];
  assign controls_counterDiff = CICC1851_controls_frameStart[25 : 18];
  always @(*) begin
    controls_twiceCompValid = CICC1851_controls_frameStart[26];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_6_HOLD : begin
      end
      controlStateMachine_enumDef_6_PASS : begin
      end
      controlStateMachine_enumDef_6_ONCE : begin
      end
      controlStateMachine_enumDef_6_TWICE : begin
        controls_twiceCompValid = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_twiceMode = CICC1851_controls_frameStart[29 : 27];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_6_HOLD : begin
      end
      controlStateMachine_enumDef_6_PASS : begin
      end
      controlStateMachine_enumDef_6_ONCE : begin
      end
      controlStateMachine_enumDef_6_TWICE : begin
        if(outReachFinalRow) begin
          if(nextRowBuffer) begin
            if(outReachRowEnd) begin
              controls_twiceMode = 3'b100;
            end else begin
              controls_twiceMode = 3'b101;
            end
          end else begin
            if(outReachRowEnd) begin
              controls_twiceMode = 3'b010;
            end else begin
              controls_twiceMode = 3'b011;
            end
          end
        end else begin
          if(nextRowBuffer) begin
            controls_twiceMode = 3'b000;
          end else begin
            controls_twiceMode = 3'b001;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    validStream_ready = (controlStream_ready && startRead);
    validStream_ready = (mainAddrOneStream_ready && startRead);
    validStream_ready = (counterAddrOneStream_ready && startRead);
    validStream_ready = (mainAddrTwoStream_ready && startRead);
    validStream_ready = (counterAddrTwoStream_ready && startRead);
  end

  assign controlStream_valid = (validStream_valid && startRead);
  assign controlStream_payload_frameStart = controls_frameStart;
  assign controlStream_payload_rowEnd = controls_rowEnd;
  assign controlStream_payload_passMode = controls_passMode;
  assign controlStream_payload_passValid = controls_passValid;
  assign controlStream_payload_onceMode = controls_onceMode;
  assign controlStream_payload_onceValid = controls_onceValid;
  assign controlStream_payload_mainCompare = controls_mainCompare;
  assign controlStream_payload_counterCompare = controls_counterCompare;
  assign controlStream_payload_mainDiff = controls_mainDiff;
  assign controlStream_payload_counterDiff = controls_counterDiff;
  assign controlStream_payload_twiceCompValid = controls_twiceCompValid;
  assign controlStream_payload_twiceMode = controls_twiceMode;
  assign mainAddrOneStream_valid = (validStream_valid && startRead);
  assign mainAddrOneStream_payload = mainAddrOne;
  assign counterAddrOneStream_valid = (validStream_valid && startRead);
  assign counterAddrOneStream_payload = counterAddrOne;
  assign mainAddrTwoStream_valid = (validStream_valid && startRead);
  assign mainAddrTwoStream_payload = mainAddrTwo;
  assign counterAddrTwoStream_valid = (validStream_valid && startRead);
  assign counterAddrTwoStream_payload = counterAddrTwo;
  assign mainAddrOneStream_ready = (! mainAddrOneStream_rValid);
  assign mainAddrOneStream_s2mPipe_valid = (mainAddrOneStream_valid || mainAddrOneStream_rValid);
  assign mainAddrOneStream_s2mPipe_payload = (mainAddrOneStream_rValid ? mainAddrOneStream_rData : mainAddrOneStream_payload);
  always @(*) begin
    mainAddrOneStream_s2mPipe_ready = mainAddrOneStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368) begin
      mainAddrOneStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368 = (! mainAddrOneStream_s2mPipe_m2sPipe_valid);
  assign mainAddrOneStream_s2mPipe_m2sPipe_valid = mainAddrOneStream_s2mPipe_rValid;
  assign mainAddrOneStream_s2mPipe_m2sPipe_payload = mainAddrOneStream_s2mPipe_rData;
  assign mainAddrOneStream_s2mPipe_m2sPipe_ready = ((! CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready) || CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready = CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_mainOnePixelStream_payload = CICC1851_lineBufferOne_port0;
  assign CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_1 = readStage_mainOnePixelStream_ready;
    if(when_Stream_l368_1) begin
      CICC1851_1 = 1'b1;
    end
  end

  assign when_Stream_l368_1 = (! readStage_mainOnePixelStream_valid);
  assign readStage_mainOnePixelStream_valid = CICC1851_readStage_mainOnePixelStream_valid;
  assign readStage_mainOnePixelStream_payload = CICC1851_readStage_mainOnePixelStream_payload_2;
  assign counterAddrOneStream_ready = (! counterAddrOneStream_rValid);
  assign counterAddrOneStream_s2mPipe_valid = (counterAddrOneStream_valid || counterAddrOneStream_rValid);
  assign counterAddrOneStream_s2mPipe_payload = (counterAddrOneStream_rValid ? counterAddrOneStream_rData : counterAddrOneStream_payload);
  always @(*) begin
    counterAddrOneStream_s2mPipe_ready = counterAddrOneStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_2) begin
      counterAddrOneStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_2 = (! counterAddrOneStream_s2mPipe_m2sPipe_valid);
  assign counterAddrOneStream_s2mPipe_m2sPipe_valid = counterAddrOneStream_s2mPipe_rValid;
  assign counterAddrOneStream_s2mPipe_m2sPipe_payload = counterAddrOneStream_s2mPipe_rData;
  assign counterAddrOneStream_s2mPipe_m2sPipe_ready = ((! CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready) || CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready = CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_counterOnePixelStream_payload = CICC1851_lineBufferOne_port1;
  assign CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_2 = readStage_counterOnePixelStream_ready;
    if(when_Stream_l368_3) begin
      CICC1851_2 = 1'b1;
    end
  end

  assign when_Stream_l368_3 = (! readStage_counterOnePixelStream_valid);
  assign readStage_counterOnePixelStream_valid = CICC1851_readStage_counterOnePixelStream_valid;
  assign readStage_counterOnePixelStream_payload = CICC1851_readStage_counterOnePixelStream_payload_2;
  assign mainAddrTwoStream_ready = (! mainAddrTwoStream_rValid);
  assign mainAddrTwoStream_s2mPipe_valid = (mainAddrTwoStream_valid || mainAddrTwoStream_rValid);
  assign mainAddrTwoStream_s2mPipe_payload = (mainAddrTwoStream_rValid ? mainAddrTwoStream_rData : mainAddrTwoStream_payload);
  always @(*) begin
    mainAddrTwoStream_s2mPipe_ready = mainAddrTwoStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_4) begin
      mainAddrTwoStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_4 = (! mainAddrTwoStream_s2mPipe_m2sPipe_valid);
  assign mainAddrTwoStream_s2mPipe_m2sPipe_valid = mainAddrTwoStream_s2mPipe_rValid;
  assign mainAddrTwoStream_s2mPipe_m2sPipe_payload = mainAddrTwoStream_s2mPipe_rData;
  assign mainAddrTwoStream_s2mPipe_m2sPipe_ready = ((! CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready) || CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready = CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_mainTwoPixelStream_payload = CICC1851_lineBufferTwo_port0;
  assign CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_3 = readStage_mainTwoPixelStream_ready;
    if(when_Stream_l368_5) begin
      CICC1851_3 = 1'b1;
    end
  end

  assign when_Stream_l368_5 = (! readStage_mainTwoPixelStream_valid);
  assign readStage_mainTwoPixelStream_valid = CICC1851_readStage_mainTwoPixelStream_valid;
  assign readStage_mainTwoPixelStream_payload = CICC1851_readStage_mainTwoPixelStream_payload_2;
  assign counterAddrTwoStream_ready = (! counterAddrTwoStream_rValid);
  assign counterAddrTwoStream_s2mPipe_valid = (counterAddrTwoStream_valid || counterAddrTwoStream_rValid);
  assign counterAddrTwoStream_s2mPipe_payload = (counterAddrTwoStream_rValid ? counterAddrTwoStream_rData : counterAddrTwoStream_payload);
  always @(*) begin
    counterAddrTwoStream_s2mPipe_ready = counterAddrTwoStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_6) begin
      counterAddrTwoStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_6 = (! counterAddrTwoStream_s2mPipe_m2sPipe_valid);
  assign counterAddrTwoStream_s2mPipe_m2sPipe_valid = counterAddrTwoStream_s2mPipe_rValid;
  assign counterAddrTwoStream_s2mPipe_m2sPipe_payload = counterAddrTwoStream_s2mPipe_rData;
  assign counterAddrTwoStream_s2mPipe_m2sPipe_ready = ((! CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready) || CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready = CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_counterTwoPixelStream_payload = CICC1851_lineBufferTwo_port1;
  assign CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_4 = readStage_counterTwoPixelStream_ready;
    if(when_Stream_l368_7) begin
      CICC1851_4 = 1'b1;
    end
  end

  assign when_Stream_l368_7 = (! readStage_counterTwoPixelStream_valid);
  assign readStage_counterTwoPixelStream_valid = CICC1851_readStage_counterTwoPixelStream_valid;
  assign readStage_counterTwoPixelStream_payload = CICC1851_readStage_counterTwoPixelStream_payload_2;
  assign controlStream_ready = (! controlStream_rValid);
  assign controlStream_s2mPipe_valid = (controlStream_valid || controlStream_rValid);
  assign controlStream_s2mPipe_payload_frameStart = (controlStream_rValid ? controlStream_rData_frameStart : controlStream_payload_frameStart);
  assign controlStream_s2mPipe_payload_rowEnd = (controlStream_rValid ? controlStream_rData_rowEnd : controlStream_payload_rowEnd);
  assign controlStream_s2mPipe_payload_passMode = (controlStream_rValid ? controlStream_rData_passMode : controlStream_payload_passMode);
  assign controlStream_s2mPipe_payload_passValid = (controlStream_rValid ? controlStream_rData_passValid : controlStream_payload_passValid);
  assign controlStream_s2mPipe_payload_onceMode = (controlStream_rValid ? controlStream_rData_onceMode : controlStream_payload_onceMode);
  assign controlStream_s2mPipe_payload_onceValid = (controlStream_rValid ? controlStream_rData_onceValid : controlStream_payload_onceValid);
  assign controlStream_s2mPipe_payload_mainCompare = (controlStream_rValid ? controlStream_rData_mainCompare : controlStream_payload_mainCompare);
  assign controlStream_s2mPipe_payload_counterCompare = (controlStream_rValid ? controlStream_rData_counterCompare : controlStream_payload_counterCompare);
  assign controlStream_s2mPipe_payload_mainDiff = (controlStream_rValid ? controlStream_rData_mainDiff : controlStream_payload_mainDiff);
  assign controlStream_s2mPipe_payload_counterDiff = (controlStream_rValid ? controlStream_rData_counterDiff : controlStream_payload_counterDiff);
  assign controlStream_s2mPipe_payload_twiceCompValid = (controlStream_rValid ? controlStream_rData_twiceCompValid : controlStream_payload_twiceCompValid);
  assign controlStream_s2mPipe_payload_twiceMode = (controlStream_rValid ? controlStream_rData_twiceMode : controlStream_payload_twiceMode);
  always @(*) begin
    controlStream_s2mPipe_ready = controlStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_8) begin
      controlStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_8 = (! controlStream_s2mPipe_m2sPipe_valid);
  assign controlStream_s2mPipe_m2sPipe_valid = controlStream_s2mPipe_rValid;
  assign controlStream_s2mPipe_m2sPipe_payload_frameStart = controlStream_s2mPipe_rData_frameStart;
  assign controlStream_s2mPipe_m2sPipe_payload_rowEnd = controlStream_s2mPipe_rData_rowEnd;
  assign controlStream_s2mPipe_m2sPipe_payload_passMode = controlStream_s2mPipe_rData_passMode;
  assign controlStream_s2mPipe_m2sPipe_payload_passValid = controlStream_s2mPipe_rData_passValid;
  assign controlStream_s2mPipe_m2sPipe_payload_onceMode = controlStream_s2mPipe_rData_onceMode;
  assign controlStream_s2mPipe_m2sPipe_payload_onceValid = controlStream_s2mPipe_rData_onceValid;
  assign controlStream_s2mPipe_m2sPipe_payload_mainCompare = controlStream_s2mPipe_rData_mainCompare;
  assign controlStream_s2mPipe_m2sPipe_payload_counterCompare = controlStream_s2mPipe_rData_counterCompare;
  assign controlStream_s2mPipe_m2sPipe_payload_mainDiff = controlStream_s2mPipe_rData_mainDiff;
  assign controlStream_s2mPipe_m2sPipe_payload_counterDiff = controlStream_s2mPipe_rData_counterDiff;
  assign controlStream_s2mPipe_m2sPipe_payload_twiceCompValid = controlStream_s2mPipe_rData_twiceCompValid;
  assign controlStream_s2mPipe_m2sPipe_payload_twiceMode = controlStream_s2mPipe_rData_twiceMode;
  always @(*) begin
    controlStream_s2mPipe_m2sPipe_ready = controlStream_s2mPipe_m2sPipe_m2sPipe_ready;
    if(when_Stream_l368_9) begin
      controlStream_s2mPipe_m2sPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_9 = (! controlStream_s2mPipe_m2sPipe_m2sPipe_valid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_valid = controlStream_s2mPipe_m2sPipe_rValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_frameStart = controlStream_s2mPipe_m2sPipe_rData_frameStart;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_rowEnd = controlStream_s2mPipe_m2sPipe_rData_rowEnd;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passMode = controlStream_s2mPipe_m2sPipe_rData_passMode;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passValid = controlStream_s2mPipe_m2sPipe_rData_passValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceMode = controlStream_s2mPipe_m2sPipe_rData_onceMode;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceValid = controlStream_s2mPipe_m2sPipe_rData_onceValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainCompare = controlStream_s2mPipe_m2sPipe_rData_mainCompare;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterCompare = controlStream_s2mPipe_m2sPipe_rData_counterCompare;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDiff = controlStream_s2mPipe_m2sPipe_rData_mainDiff;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDiff = controlStream_s2mPipe_m2sPipe_rData_counterDiff;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceCompValid = controlStream_s2mPipe_m2sPipe_rData_twiceCompValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceMode = controlStream_s2mPipe_m2sPipe_rData_twiceMode;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_ready = (! controlStream_s2mPipe_m2sPipe_m2sPipe_rValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_valid = (controlStream_s2mPipe_m2sPipe_m2sPipe_valid || controlStream_s2mPipe_m2sPipe_m2sPipe_rValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_frameStart = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_frameStart : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_frameStart);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_rowEnd = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_rowEnd : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_rowEnd);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_passMode = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_passMode : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passMode);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_passValid = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_passValid : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_onceMode = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_onceMode : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceMode);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_onceValid = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_onceValid : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainCompare = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainCompare : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainCompare);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterCompare = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterCompare : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterCompare);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainDiff = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainDiff : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDiff);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterDiff = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterDiff : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDiff);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_twiceCompValid = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_twiceCompValid : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceCompValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_twiceMode = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_twiceMode : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceMode);
  always @(*) begin
    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready = readStage_controlPipe_ready;
    if(when_Stream_l368_10) begin
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_10 = (! readStage_controlPipe_valid);
  assign readStage_controlPipe_valid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rValid;
  assign readStage_controlPipe_payload_frameStart = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_frameStart;
  assign readStage_controlPipe_payload_rowEnd = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_rowEnd;
  assign readStage_controlPipe_payload_passMode = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_passMode;
  assign readStage_controlPipe_payload_passValid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_passValid;
  assign readStage_controlPipe_payload_onceMode = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_onceMode;
  assign readStage_controlPipe_payload_onceValid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_onceValid;
  assign readStage_controlPipe_payload_mainCompare = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainCompare;
  assign readStage_controlPipe_payload_counterCompare = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterCompare;
  assign readStage_controlPipe_payload_mainDiff = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainDiff;
  assign readStage_controlPipe_payload_counterDiff = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterDiff;
  assign readStage_controlPipe_payload_twiceCompValid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_twiceCompValid;
  assign readStage_controlPipe_payload_twiceMode = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_twiceMode;
  assign readStage_mainOnePixelStream_ready = (! readStage_mainOnePixelStream_rValid);
  assign readStage_mainOnePixelStream_s2mPipe_valid = (readStage_mainOnePixelStream_valid || readStage_mainOnePixelStream_rValid);
  assign readStage_mainOnePixelStream_s2mPipe_payload = (readStage_mainOnePixelStream_rValid ? readStage_mainOnePixelStream_rData : readStage_mainOnePixelStream_payload);
  always @(*) begin
    readStage_mainOnePixelStream_s2mPipe_ready = compareStage_mainOnePixelStream_ready;
    if(when_Stream_l368_11) begin
      readStage_mainOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_11 = (! compareStage_mainOnePixelStream_valid);
  assign compareStage_mainOnePixelStream_valid = readStage_mainOnePixelStream_s2mPipe_rValid;
  assign compareStage_mainOnePixelStream_payload = readStage_mainOnePixelStream_s2mPipe_rData;
  assign readStage_counterOnePixelStream_ready = (! readStage_counterOnePixelStream_rValid);
  assign readStage_counterOnePixelStream_s2mPipe_valid = (readStage_counterOnePixelStream_valid || readStage_counterOnePixelStream_rValid);
  assign readStage_counterOnePixelStream_s2mPipe_payload = (readStage_counterOnePixelStream_rValid ? readStage_counterOnePixelStream_rData : readStage_counterOnePixelStream_payload);
  always @(*) begin
    readStage_counterOnePixelStream_s2mPipe_ready = compareStage_counterOnePixelStream_ready;
    if(when_Stream_l368_12) begin
      readStage_counterOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_12 = (! compareStage_counterOnePixelStream_valid);
  assign compareStage_counterOnePixelStream_valid = readStage_counterOnePixelStream_s2mPipe_rValid;
  assign compareStage_counterOnePixelStream_payload = readStage_counterOnePixelStream_s2mPipe_rData;
  assign readStage_mainTwoPixelStream_ready = (! readStage_mainTwoPixelStream_rValid);
  assign readStage_mainTwoPixelStream_s2mPipe_valid = (readStage_mainTwoPixelStream_valid || readStage_mainTwoPixelStream_rValid);
  assign readStage_mainTwoPixelStream_s2mPipe_payload = (readStage_mainTwoPixelStream_rValid ? readStage_mainTwoPixelStream_rData : readStage_mainTwoPixelStream_payload);
  always @(*) begin
    readStage_mainTwoPixelStream_s2mPipe_ready = compareStage_mainTwoPixelStream_ready;
    if(when_Stream_l368_13) begin
      readStage_mainTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_13 = (! compareStage_mainTwoPixelStream_valid);
  assign compareStage_mainTwoPixelStream_valid = readStage_mainTwoPixelStream_s2mPipe_rValid;
  assign compareStage_mainTwoPixelStream_payload = readStage_mainTwoPixelStream_s2mPipe_rData;
  assign readStage_counterTwoPixelStream_ready = (! readStage_counterTwoPixelStream_rValid);
  assign readStage_counterTwoPixelStream_s2mPipe_valid = (readStage_counterTwoPixelStream_valid || readStage_counterTwoPixelStream_rValid);
  assign readStage_counterTwoPixelStream_s2mPipe_payload = (readStage_counterTwoPixelStream_rValid ? readStage_counterTwoPixelStream_rData : readStage_counterTwoPixelStream_payload);
  always @(*) begin
    readStage_counterTwoPixelStream_s2mPipe_ready = compareStage_counterTwoPixelStream_ready;
    if(when_Stream_l368_14) begin
      readStage_counterTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_14 = (! compareStage_counterTwoPixelStream_valid);
  assign compareStage_counterTwoPixelStream_valid = readStage_counterTwoPixelStream_s2mPipe_rValid;
  assign compareStage_counterTwoPixelStream_payload = readStage_counterTwoPixelStream_s2mPipe_rData;
  always @(*) begin
    CICC1851_readStage_controlPipe_translated_payload_mainCompare = readStage_controlPipe_payload_mainCompare;
    if(readStage_controlPipe_payload_onceValid) begin
      case(readStage_controlPipe_payload_onceMode)
        3'b000 : begin
          if(when_SuperResolutionPart1_l205) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        3'b001 : begin
          if(when_SuperResolutionPart1_l209) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        3'b010 : begin
          if(when_SuperResolutionPart1_l213) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        3'b011 : begin
          if(when_SuperResolutionPart1_l217) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        3'b100 : begin
          CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
        end
        3'b101 : begin
          CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
        end
        default : begin
        end
      endcase
    end
    if(readStage_controlPipe_payload_twiceCompValid) begin
      case(readStage_controlPipe_payload_twiceMode)
        3'b000 : begin
          if(when_SuperResolutionPart1_l228) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        3'b001 : begin
          if(when_SuperResolutionPart1_l234) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        3'b010 : begin
          CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
        end
        3'b011 : begin
          if(when_SuperResolutionPart1_l241) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        3'b100 : begin
          CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
        end
        3'b101 : begin
          if(when_SuperResolutionPart1_l246) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    CICC1851_readStage_controlPipe_translated_payload_counterCompare = readStage_controlPipe_payload_counterCompare;
    if(readStage_controlPipe_payload_twiceCompValid) begin
      case(readStage_controlPipe_payload_twiceMode)
        3'b000 : begin
          if(when_SuperResolutionPart1_l230) begin
            CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
          end
        end
        3'b001 : begin
          if(when_SuperResolutionPart1_l236) begin
            CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
          end
        end
        default : begin
        end
      endcase
    end
  end

  assign when_SuperResolutionPart1_l205 = (readStage_counterOnePixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart1_l209 = (readStage_counterTwoPixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart1_l213 = (readStage_mainTwoPixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart1_l217 = (readStage_mainOnePixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart1_l228 = (readStage_mainTwoPixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart1_l230 = (readStage_counterOnePixelStream_payload <= readStage_counterTwoPixelStream_payload);
  assign when_SuperResolutionPart1_l234 = (readStage_mainOnePixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart1_l236 = (readStage_counterTwoPixelStream_payload <= readStage_counterOnePixelStream_payload);
  assign when_SuperResolutionPart1_l241 = (readStage_counterTwoPixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart1_l246 = (readStage_counterOnePixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign readStage_controlPipe_translated_valid = readStage_controlPipe_valid;
  assign readStage_controlPipe_ready = readStage_controlPipe_translated_ready;
  assign readStage_controlPipe_translated_payload_frameStart = readStage_controlPipe_payload_frameStart;
  assign readStage_controlPipe_translated_payload_rowEnd = readStage_controlPipe_payload_rowEnd;
  assign readStage_controlPipe_translated_payload_passMode = readStage_controlPipe_payload_passMode;
  assign readStage_controlPipe_translated_payload_passValid = readStage_controlPipe_payload_passValid;
  assign readStage_controlPipe_translated_payload_onceMode = readStage_controlPipe_payload_onceMode;
  assign readStage_controlPipe_translated_payload_onceValid = readStage_controlPipe_payload_onceValid;
  assign readStage_controlPipe_translated_payload_mainCompare = CICC1851_readStage_controlPipe_translated_payload_mainCompare;
  assign readStage_controlPipe_translated_payload_counterCompare = CICC1851_readStage_controlPipe_translated_payload_counterCompare;
  assign readStage_controlPipe_translated_payload_mainDiff = readStage_controlPipe_payload_mainDiff;
  assign readStage_controlPipe_translated_payload_counterDiff = readStage_controlPipe_payload_counterDiff;
  assign readStage_controlPipe_translated_payload_twiceCompValid = readStage_controlPipe_payload_twiceCompValid;
  assign readStage_controlPipe_translated_payload_twiceMode = readStage_controlPipe_payload_twiceMode;
  assign readStage_controlPipe_translated_ready = (! readStage_controlPipe_translated_rValid);
  assign readStage_controlPipe_translated_s2mPipe_valid = (readStage_controlPipe_translated_valid || readStage_controlPipe_translated_rValid);
  assign readStage_controlPipe_translated_s2mPipe_payload_frameStart = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_frameStart : readStage_controlPipe_translated_payload_frameStart);
  assign readStage_controlPipe_translated_s2mPipe_payload_rowEnd = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_rowEnd : readStage_controlPipe_translated_payload_rowEnd);
  assign readStage_controlPipe_translated_s2mPipe_payload_passMode = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_passMode : readStage_controlPipe_translated_payload_passMode);
  assign readStage_controlPipe_translated_s2mPipe_payload_passValid = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_passValid : readStage_controlPipe_translated_payload_passValid);
  assign readStage_controlPipe_translated_s2mPipe_payload_onceMode = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_onceMode : readStage_controlPipe_translated_payload_onceMode);
  assign readStage_controlPipe_translated_s2mPipe_payload_onceValid = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_onceValid : readStage_controlPipe_translated_payload_onceValid);
  assign readStage_controlPipe_translated_s2mPipe_payload_mainCompare = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_mainCompare : readStage_controlPipe_translated_payload_mainCompare);
  assign readStage_controlPipe_translated_s2mPipe_payload_counterCompare = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_counterCompare : readStage_controlPipe_translated_payload_counterCompare);
  assign readStage_controlPipe_translated_s2mPipe_payload_mainDiff = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_mainDiff : readStage_controlPipe_translated_payload_mainDiff);
  assign readStage_controlPipe_translated_s2mPipe_payload_counterDiff = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_counterDiff : readStage_controlPipe_translated_payload_counterDiff);
  assign readStage_controlPipe_translated_s2mPipe_payload_twiceCompValid = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_twiceCompValid : readStage_controlPipe_translated_payload_twiceCompValid);
  assign readStage_controlPipe_translated_s2mPipe_payload_twiceMode = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_twiceMode : readStage_controlPipe_translated_payload_twiceMode);
  always @(*) begin
    readStage_controlPipe_translated_s2mPipe_ready = compareStage_controlPipe_ready;
    if(when_Stream_l368_15) begin
      readStage_controlPipe_translated_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_15 = (! compareStage_controlPipe_valid);
  assign compareStage_controlPipe_valid = readStage_controlPipe_translated_s2mPipe_rValid;
  assign compareStage_controlPipe_payload_frameStart = readStage_controlPipe_translated_s2mPipe_rData_frameStart;
  assign compareStage_controlPipe_payload_rowEnd = readStage_controlPipe_translated_s2mPipe_rData_rowEnd;
  assign compareStage_controlPipe_payload_passMode = readStage_controlPipe_translated_s2mPipe_rData_passMode;
  assign compareStage_controlPipe_payload_passValid = readStage_controlPipe_translated_s2mPipe_rData_passValid;
  assign compareStage_controlPipe_payload_onceMode = readStage_controlPipe_translated_s2mPipe_rData_onceMode;
  assign compareStage_controlPipe_payload_onceValid = readStage_controlPipe_translated_s2mPipe_rData_onceValid;
  assign compareStage_controlPipe_payload_mainCompare = readStage_controlPipe_translated_s2mPipe_rData_mainCompare;
  assign compareStage_controlPipe_payload_counterCompare = readStage_controlPipe_translated_s2mPipe_rData_counterCompare;
  assign compareStage_controlPipe_payload_mainDiff = readStage_controlPipe_translated_s2mPipe_rData_mainDiff;
  assign compareStage_controlPipe_payload_counterDiff = readStage_controlPipe_translated_s2mPipe_rData_counterDiff;
  assign compareStage_controlPipe_payload_twiceCompValid = readStage_controlPipe_translated_s2mPipe_rData_twiceCompValid;
  assign compareStage_controlPipe_payload_twiceMode = readStage_controlPipe_translated_s2mPipe_rData_twiceMode;
  assign compareStage_mainOnePixelStream_ready = (! compareStage_mainOnePixelStream_rValid);
  assign compareStage_mainOnePixelStream_s2mPipe_valid = (compareStage_mainOnePixelStream_valid || compareStage_mainOnePixelStream_rValid);
  assign compareStage_mainOnePixelStream_s2mPipe_payload = (compareStage_mainOnePixelStream_rValid ? compareStage_mainOnePixelStream_rData : compareStage_mainOnePixelStream_payload);
  always @(*) begin
    compareStage_mainOnePixelStream_s2mPipe_ready = diffStage_mainOnePixelStream_ready;
    if(when_Stream_l368_16) begin
      compareStage_mainOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_16 = (! diffStage_mainOnePixelStream_valid);
  assign diffStage_mainOnePixelStream_valid = compareStage_mainOnePixelStream_s2mPipe_rValid;
  assign diffStage_mainOnePixelStream_payload = compareStage_mainOnePixelStream_s2mPipe_rData;
  assign compareStage_counterOnePixelStream_ready = (! compareStage_counterOnePixelStream_rValid);
  assign compareStage_counterOnePixelStream_s2mPipe_valid = (compareStage_counterOnePixelStream_valid || compareStage_counterOnePixelStream_rValid);
  assign compareStage_counterOnePixelStream_s2mPipe_payload = (compareStage_counterOnePixelStream_rValid ? compareStage_counterOnePixelStream_rData : compareStage_counterOnePixelStream_payload);
  always @(*) begin
    compareStage_counterOnePixelStream_s2mPipe_ready = diffStage_counterOnePixelStream_ready;
    if(when_Stream_l368_17) begin
      compareStage_counterOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_17 = (! diffStage_counterOnePixelStream_valid);
  assign diffStage_counterOnePixelStream_valid = compareStage_counterOnePixelStream_s2mPipe_rValid;
  assign diffStage_counterOnePixelStream_payload = compareStage_counterOnePixelStream_s2mPipe_rData;
  assign compareStage_mainTwoPixelStream_ready = (! compareStage_mainTwoPixelStream_rValid);
  assign compareStage_mainTwoPixelStream_s2mPipe_valid = (compareStage_mainTwoPixelStream_valid || compareStage_mainTwoPixelStream_rValid);
  assign compareStage_mainTwoPixelStream_s2mPipe_payload = (compareStage_mainTwoPixelStream_rValid ? compareStage_mainTwoPixelStream_rData : compareStage_mainTwoPixelStream_payload);
  always @(*) begin
    compareStage_mainTwoPixelStream_s2mPipe_ready = diffStage_mainTwoPixelStream_ready;
    if(when_Stream_l368_18) begin
      compareStage_mainTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_18 = (! diffStage_mainTwoPixelStream_valid);
  assign diffStage_mainTwoPixelStream_valid = compareStage_mainTwoPixelStream_s2mPipe_rValid;
  assign diffStage_mainTwoPixelStream_payload = compareStage_mainTwoPixelStream_s2mPipe_rData;
  assign compareStage_counterTwoPixelStream_ready = (! compareStage_counterTwoPixelStream_rValid);
  assign compareStage_counterTwoPixelStream_s2mPipe_valid = (compareStage_counterTwoPixelStream_valid || compareStage_counterTwoPixelStream_rValid);
  assign compareStage_counterTwoPixelStream_s2mPipe_payload = (compareStage_counterTwoPixelStream_rValid ? compareStage_counterTwoPixelStream_rData : compareStage_counterTwoPixelStream_payload);
  always @(*) begin
    compareStage_counterTwoPixelStream_s2mPipe_ready = diffStage_counterTwoPixelStream_ready;
    if(when_Stream_l368_19) begin
      compareStage_counterTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_19 = (! diffStage_counterTwoPixelStream_valid);
  assign diffStage_counterTwoPixelStream_valid = compareStage_counterTwoPixelStream_s2mPipe_rValid;
  assign diffStage_counterTwoPixelStream_payload = compareStage_counterTwoPixelStream_s2mPipe_rData;
  always @(*) begin
    CICC1851_compareStage_controlPipe_translated_payload_mainDiff = compareStage_controlPipe_payload_mainDiff;
    if(compareStage_controlPipe_payload_onceValid) begin
      case(compareStage_controlPipe_payload_onceMode)
        3'b000 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_counterOnePixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterOnePixelStream_payload - compareStage_mainOnePixelStream_payload);
          end
        end
        3'b001 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterTwoPixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainTwoPixelStream_payload);
          end
        end
        3'b010 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_mainTwoPixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_mainOnePixelStream_payload);
          end
        end
        3'b011 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_mainOnePixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_mainTwoPixelStream_payload);
          end
        end
        3'b100 : begin
          CICC1851_compareStage_controlPipe_translated_payload_mainDiff = 8'h0;
        end
        3'b101 : begin
          CICC1851_compareStage_controlPipe_translated_payload_mainDiff = 8'h0;
        end
        default : begin
        end
      endcase
    end
    if(compareStage_controlPipe_payload_twiceCompValid) begin
      case(compareStage_controlPipe_payload_twiceMode)
        3'b000 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_mainTwoPixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_mainOnePixelStream_payload);
          end
        end
        3'b001 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_mainOnePixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_mainTwoPixelStream_payload);
          end
        end
        3'b010 : begin
          CICC1851_compareStage_controlPipe_translated_payload_mainDiff = 8'h0;
        end
        3'b011 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterTwoPixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainTwoPixelStream_payload);
          end
        end
        3'b100 : begin
          CICC1851_compareStage_controlPipe_translated_payload_mainDiff = 8'h0;
        end
        3'b101 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_counterOnePixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterOnePixelStream_payload - compareStage_mainOnePixelStream_payload);
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    CICC1851_compareStage_controlPipe_translated_payload_counterDiff = compareStage_controlPipe_payload_counterDiff;
    if(compareStage_controlPipe_payload_twiceCompValid) begin
      case(compareStage_controlPipe_payload_twiceMode)
        3'b000 : begin
          if(compareStage_controlPipe_payload_counterCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterTwoPixelStream_payload - compareStage_counterOnePixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterOnePixelStream_payload - compareStage_counterTwoPixelStream_payload);
          end
        end
        3'b001 : begin
          if(compareStage_controlPipe_payload_counterCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterOnePixelStream_payload - compareStage_counterTwoPixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterTwoPixelStream_payload - compareStage_counterOnePixelStream_payload);
          end
        end
        default : begin
        end
      endcase
    end
  end

  assign compareStage_controlPipe_translated_valid = compareStage_controlPipe_valid;
  assign compareStage_controlPipe_ready = compareStage_controlPipe_translated_ready;
  assign compareStage_controlPipe_translated_payload_frameStart = compareStage_controlPipe_payload_frameStart;
  assign compareStage_controlPipe_translated_payload_rowEnd = compareStage_controlPipe_payload_rowEnd;
  assign compareStage_controlPipe_translated_payload_passMode = compareStage_controlPipe_payload_passMode;
  assign compareStage_controlPipe_translated_payload_passValid = compareStage_controlPipe_payload_passValid;
  assign compareStage_controlPipe_translated_payload_onceMode = compareStage_controlPipe_payload_onceMode;
  assign compareStage_controlPipe_translated_payload_onceValid = compareStage_controlPipe_payload_onceValid;
  assign compareStage_controlPipe_translated_payload_mainCompare = compareStage_controlPipe_payload_mainCompare;
  assign compareStage_controlPipe_translated_payload_counterCompare = compareStage_controlPipe_payload_counterCompare;
  assign compareStage_controlPipe_translated_payload_mainDiff = CICC1851_compareStage_controlPipe_translated_payload_mainDiff;
  assign compareStage_controlPipe_translated_payload_counterDiff = CICC1851_compareStage_controlPipe_translated_payload_counterDiff;
  assign compareStage_controlPipe_translated_payload_twiceCompValid = compareStage_controlPipe_payload_twiceCompValid;
  assign compareStage_controlPipe_translated_payload_twiceMode = compareStage_controlPipe_payload_twiceMode;
  assign compareStage_controlPipe_translated_ready = (! compareStage_controlPipe_translated_rValid);
  assign compareStage_controlPipe_translated_s2mPipe_valid = (compareStage_controlPipe_translated_valid || compareStage_controlPipe_translated_rValid);
  assign compareStage_controlPipe_translated_s2mPipe_payload_frameStart = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_frameStart : compareStage_controlPipe_translated_payload_frameStart);
  assign compareStage_controlPipe_translated_s2mPipe_payload_rowEnd = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_rowEnd : compareStage_controlPipe_translated_payload_rowEnd);
  assign compareStage_controlPipe_translated_s2mPipe_payload_passMode = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_passMode : compareStage_controlPipe_translated_payload_passMode);
  assign compareStage_controlPipe_translated_s2mPipe_payload_passValid = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_passValid : compareStage_controlPipe_translated_payload_passValid);
  assign compareStage_controlPipe_translated_s2mPipe_payload_onceMode = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_onceMode : compareStage_controlPipe_translated_payload_onceMode);
  assign compareStage_controlPipe_translated_s2mPipe_payload_onceValid = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_onceValid : compareStage_controlPipe_translated_payload_onceValid);
  assign compareStage_controlPipe_translated_s2mPipe_payload_mainCompare = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_mainCompare : compareStage_controlPipe_translated_payload_mainCompare);
  assign compareStage_controlPipe_translated_s2mPipe_payload_counterCompare = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_counterCompare : compareStage_controlPipe_translated_payload_counterCompare);
  assign compareStage_controlPipe_translated_s2mPipe_payload_mainDiff = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_mainDiff : compareStage_controlPipe_translated_payload_mainDiff);
  assign compareStage_controlPipe_translated_s2mPipe_payload_counterDiff = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_counterDiff : compareStage_controlPipe_translated_payload_counterDiff);
  assign compareStage_controlPipe_translated_s2mPipe_payload_twiceCompValid = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_twiceCompValid : compareStage_controlPipe_translated_payload_twiceCompValid);
  assign compareStage_controlPipe_translated_s2mPipe_payload_twiceMode = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_twiceMode : compareStage_controlPipe_translated_payload_twiceMode);
  always @(*) begin
    compareStage_controlPipe_translated_s2mPipe_ready = diffStage_controlPipe_ready;
    if(when_Stream_l368_20) begin
      compareStage_controlPipe_translated_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_20 = (! diffStage_controlPipe_valid);
  assign diffStage_controlPipe_valid = compareStage_controlPipe_translated_s2mPipe_rValid;
  assign diffStage_controlPipe_payload_frameStart = compareStage_controlPipe_translated_s2mPipe_rData_frameStart;
  assign diffStage_controlPipe_payload_rowEnd = compareStage_controlPipe_translated_s2mPipe_rData_rowEnd;
  assign diffStage_controlPipe_payload_passMode = compareStage_controlPipe_translated_s2mPipe_rData_passMode;
  assign diffStage_controlPipe_payload_passValid = compareStage_controlPipe_translated_s2mPipe_rData_passValid;
  assign diffStage_controlPipe_payload_onceMode = compareStage_controlPipe_translated_s2mPipe_rData_onceMode;
  assign diffStage_controlPipe_payload_onceValid = compareStage_controlPipe_translated_s2mPipe_rData_onceValid;
  assign diffStage_controlPipe_payload_mainCompare = compareStage_controlPipe_translated_s2mPipe_rData_mainCompare;
  assign diffStage_controlPipe_payload_counterCompare = compareStage_controlPipe_translated_s2mPipe_rData_counterCompare;
  assign diffStage_controlPipe_payload_mainDiff = compareStage_controlPipe_translated_s2mPipe_rData_mainDiff;
  assign diffStage_controlPipe_payload_counterDiff = compareStage_controlPipe_translated_s2mPipe_rData_counterDiff;
  assign diffStage_controlPipe_payload_twiceCompValid = compareStage_controlPipe_translated_s2mPipe_rData_twiceCompValid;
  assign diffStage_controlPipe_payload_twiceMode = compareStage_controlPipe_translated_s2mPipe_rData_twiceMode;
  assign diffStage_mainOnePixelStream_ready = (! diffStage_mainOnePixelStream_rValid);
  assign diffStage_mainOnePixelStream_s2mPipe_valid = (diffStage_mainOnePixelStream_valid || diffStage_mainOnePixelStream_rValid);
  assign diffStage_mainOnePixelStream_s2mPipe_payload = (diffStage_mainOnePixelStream_rValid ? diffStage_mainOnePixelStream_rData : diffStage_mainOnePixelStream_payload);
  always @(*) begin
    diffStage_mainOnePixelStream_s2mPipe_ready = resultStage_mainOnePixelStream_ready;
    if(when_Stream_l368_21) begin
      diffStage_mainOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_21 = (! resultStage_mainOnePixelStream_valid);
  assign resultStage_mainOnePixelStream_valid = diffStage_mainOnePixelStream_s2mPipe_rValid;
  assign resultStage_mainOnePixelStream_payload = diffStage_mainOnePixelStream_s2mPipe_rData;
  assign diffStage_counterOnePixelStream_ready = (! diffStage_counterOnePixelStream_rValid);
  assign diffStage_counterOnePixelStream_s2mPipe_valid = (diffStage_counterOnePixelStream_valid || diffStage_counterOnePixelStream_rValid);
  assign diffStage_counterOnePixelStream_s2mPipe_payload = (diffStage_counterOnePixelStream_rValid ? diffStage_counterOnePixelStream_rData : diffStage_counterOnePixelStream_payload);
  always @(*) begin
    diffStage_counterOnePixelStream_s2mPipe_ready = resultStage_counterOnePixelStream_ready;
    if(when_Stream_l368_22) begin
      diffStage_counterOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_22 = (! resultStage_counterOnePixelStream_valid);
  assign resultStage_counterOnePixelStream_valid = diffStage_counterOnePixelStream_s2mPipe_rValid;
  assign resultStage_counterOnePixelStream_payload = diffStage_counterOnePixelStream_s2mPipe_rData;
  assign diffStage_mainTwoPixelStream_ready = (! diffStage_mainTwoPixelStream_rValid);
  assign diffStage_mainTwoPixelStream_s2mPipe_valid = (diffStage_mainTwoPixelStream_valid || diffStage_mainTwoPixelStream_rValid);
  assign diffStage_mainTwoPixelStream_s2mPipe_payload = (diffStage_mainTwoPixelStream_rValid ? diffStage_mainTwoPixelStream_rData : diffStage_mainTwoPixelStream_payload);
  always @(*) begin
    diffStage_mainTwoPixelStream_s2mPipe_ready = resultStage_mainTwoPixelStream_ready;
    if(when_Stream_l368_23) begin
      diffStage_mainTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_23 = (! resultStage_mainTwoPixelStream_valid);
  assign resultStage_mainTwoPixelStream_valid = diffStage_mainTwoPixelStream_s2mPipe_rValid;
  assign resultStage_mainTwoPixelStream_payload = diffStage_mainTwoPixelStream_s2mPipe_rData;
  assign diffStage_counterTwoPixelStream_ready = (! diffStage_counterTwoPixelStream_rValid);
  assign diffStage_counterTwoPixelStream_s2mPipe_valid = (diffStage_counterTwoPixelStream_valid || diffStage_counterTwoPixelStream_rValid);
  assign diffStage_counterTwoPixelStream_s2mPipe_payload = (diffStage_counterTwoPixelStream_rValid ? diffStage_counterTwoPixelStream_rData : diffStage_counterTwoPixelStream_payload);
  always @(*) begin
    diffStage_counterTwoPixelStream_s2mPipe_ready = resultStage_counterTwoPixelStream_ready;
    if(when_Stream_l368_24) begin
      diffStage_counterTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_24 = (! resultStage_counterTwoPixelStream_valid);
  assign resultStage_counterTwoPixelStream_valid = diffStage_counterTwoPixelStream_s2mPipe_rValid;
  assign resultStage_counterTwoPixelStream_payload = diffStage_counterTwoPixelStream_s2mPipe_rData;
  assign diffStage_controlPipe_ready = diffStage_controlPipe_fork_io_input_ready;
  assign diffStage_controlPipe_fork_io_outputs_0_ready = (! diffStage_controlPipe_fork_io_outputs_0_rValid);
  assign diffStage_controlPipe_fork_io_outputs_0_s2mPipe_valid = (diffStage_controlPipe_fork_io_outputs_0_valid || diffStage_controlPipe_fork_io_outputs_0_rValid);
  assign diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_frameStart = (diffStage_controlPipe_fork_io_outputs_0_rValid ? diffStage_controlPipe_fork_io_outputs_0_rData_frameStart : diffStage_controlPipe_fork_io_outputs_0_payload_frameStart);
  assign diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_rowEnd = (diffStage_controlPipe_fork_io_outputs_0_rValid ? diffStage_controlPipe_fork_io_outputs_0_rData_rowEnd : diffStage_controlPipe_fork_io_outputs_0_payload_rowEnd);
  assign diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_passMode = (diffStage_controlPipe_fork_io_outputs_0_rValid ? diffStage_controlPipe_fork_io_outputs_0_rData_passMode : diffStage_controlPipe_fork_io_outputs_0_payload_passMode);
  assign diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_passValid = (diffStage_controlPipe_fork_io_outputs_0_rValid ? diffStage_controlPipe_fork_io_outputs_0_rData_passValid : diffStage_controlPipe_fork_io_outputs_0_payload_passValid);
  assign diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_onceMode = (diffStage_controlPipe_fork_io_outputs_0_rValid ? diffStage_controlPipe_fork_io_outputs_0_rData_onceMode : diffStage_controlPipe_fork_io_outputs_0_payload_onceMode);
  assign diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_onceValid = (diffStage_controlPipe_fork_io_outputs_0_rValid ? diffStage_controlPipe_fork_io_outputs_0_rData_onceValid : diffStage_controlPipe_fork_io_outputs_0_payload_onceValid);
  assign diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_mainCompare = (diffStage_controlPipe_fork_io_outputs_0_rValid ? diffStage_controlPipe_fork_io_outputs_0_rData_mainCompare : diffStage_controlPipe_fork_io_outputs_0_payload_mainCompare);
  assign diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_counterCompare = (diffStage_controlPipe_fork_io_outputs_0_rValid ? diffStage_controlPipe_fork_io_outputs_0_rData_counterCompare : diffStage_controlPipe_fork_io_outputs_0_payload_counterCompare);
  assign diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_mainDiff = (diffStage_controlPipe_fork_io_outputs_0_rValid ? diffStage_controlPipe_fork_io_outputs_0_rData_mainDiff : diffStage_controlPipe_fork_io_outputs_0_payload_mainDiff);
  assign diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_counterDiff = (diffStage_controlPipe_fork_io_outputs_0_rValid ? diffStage_controlPipe_fork_io_outputs_0_rData_counterDiff : diffStage_controlPipe_fork_io_outputs_0_payload_counterDiff);
  assign diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_twiceCompValid = (diffStage_controlPipe_fork_io_outputs_0_rValid ? diffStage_controlPipe_fork_io_outputs_0_rData_twiceCompValid : diffStage_controlPipe_fork_io_outputs_0_payload_twiceCompValid);
  assign diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_twiceMode = (diffStage_controlPipe_fork_io_outputs_0_rValid ? diffStage_controlPipe_fork_io_outputs_0_rData_twiceMode : diffStage_controlPipe_fork_io_outputs_0_payload_twiceMode);
  always @(*) begin
    diffStage_controlPipe_fork_io_outputs_0_s2mPipe_ready = resultStage_controlPipe_ready;
    if(when_Stream_l368_25) begin
      diffStage_controlPipe_fork_io_outputs_0_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_25 = (! resultStage_controlPipe_valid);
  assign resultStage_controlPipe_valid = diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rValid;
  assign resultStage_controlPipe_payload_frameStart = diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_frameStart;
  assign resultStage_controlPipe_payload_rowEnd = diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_rowEnd;
  assign resultStage_controlPipe_payload_passMode = diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_passMode;
  assign resultStage_controlPipe_payload_passValid = diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_passValid;
  assign resultStage_controlPipe_payload_onceMode = diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_onceMode;
  assign resultStage_controlPipe_payload_onceValid = diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_onceValid;
  assign resultStage_controlPipe_payload_mainCompare = diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_mainCompare;
  assign resultStage_controlPipe_payload_counterCompare = diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_counterCompare;
  assign resultStage_controlPipe_payload_mainDiff = diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_mainDiff;
  assign resultStage_controlPipe_payload_counterDiff = diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_counterDiff;
  assign resultStage_controlPipe_payload_twiceCompValid = diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_twiceCompValid;
  assign resultStage_controlPipe_payload_twiceMode = diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_twiceMode;
  assign resultStage_pixelStream_valid = diffStage_controlPipe_fork_io_outputs_1_valid;
  always @(*) begin
    resultStage_pixelStream_payload = 8'h0;
    if(diffStage_controlPipe_fork_io_outputs_1_payload_passValid) begin
      if(diffStage_controlPipe_fork_io_outputs_1_payload_passMode) begin
        resultStage_pixelStream_payload = diffStage_mainTwoPixelStream_payload;
      end else begin
        resultStage_pixelStream_payload = diffStage_mainOnePixelStream_payload;
      end
    end
    if(diffStage_controlPipe_fork_io_outputs_1_payload_onceValid) begin
      case(diffStage_controlPipe_fork_io_outputs_1_payload_onceMode)
        3'b000 : begin
          if(when_SuperResolutionPart1_l339) begin
            resultStage_pixelStream_payload = diffStage_mainOnePixelStream_payload;
          end else begin
            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload[7:0];
          end
        end
        3'b001 : begin
          if(when_SuperResolutionPart1_l343) begin
            resultStage_pixelStream_payload = diffStage_mainTwoPixelStream_payload;
          end else begin
            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_2[7:0];
          end
        end
        3'b010 : begin
          if(when_SuperResolutionPart1_l347) begin
            resultStage_pixelStream_payload = diffStage_mainOnePixelStream_payload;
          end else begin
            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_4[7:0];
          end
        end
        3'b011 : begin
          if(when_SuperResolutionPart1_l351) begin
            resultStage_pixelStream_payload = diffStage_mainTwoPixelStream_payload;
          end else begin
            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_6[7:0];
          end
        end
        3'b100 : begin
          resultStage_pixelStream_payload = diffStage_mainTwoPixelStream_payload;
        end
        3'b101 : begin
          resultStage_pixelStream_payload = diffStage_mainOnePixelStream_payload;
        end
        default : begin
        end
      endcase
    end
    if(diffStage_controlPipe_fork_io_outputs_1_payload_twiceCompValid) begin
      case(diffStage_controlPipe_fork_io_outputs_1_payload_twiceMode)
        3'b000 : begin
          if(when_SuperResolutionPart1_l362) begin
            if(when_SuperResolutionPart1_l363) begin
              resultStage_pixelStream_payload = diffStage_mainOnePixelStream_payload;
            end else begin
              resultStage_pixelStream_payload = diffStage_counterTwoPixelStream_payload;
            end
          end else begin
            if(when_SuperResolutionPart1_l366) begin
              resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_8[7:0];
            end else begin
              resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_10[7:0];
            end
          end
        end
        3'b001 : begin
          if(when_SuperResolutionPart1_l371) begin
            if(when_SuperResolutionPart1_l372) begin
              resultStage_pixelStream_payload = diffStage_mainTwoPixelStream_payload;
            end else begin
              resultStage_pixelStream_payload = diffStage_counterOnePixelStream_payload;
            end
          end else begin
            if(when_SuperResolutionPart1_l375) begin
              resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_12[7:0];
            end else begin
              resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_14[7:0];
            end
          end
        end
        3'b010 : begin
          resultStage_pixelStream_payload = diffStage_mainTwoPixelStream_payload;
        end
        3'b011 : begin
          if(when_SuperResolutionPart1_l381) begin
            resultStage_pixelStream_payload = diffStage_mainTwoPixelStream_payload;
          end else begin
            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_16[7:0];
          end
        end
        3'b100 : begin
          resultStage_pixelStream_payload = diffStage_mainOnePixelStream_payload;
        end
        3'b101 : begin
          if(when_SuperResolutionPart1_l386) begin
            resultStage_pixelStream_payload = diffStage_mainOnePixelStream_payload;
          end else begin
            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_18[7:0];
          end
        end
        default : begin
        end
      endcase
    end
  end

  assign when_SuperResolutionPart1_l339 = (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart1_l343 = (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart1_l347 = (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart1_l351 = (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart1_l362 = ((inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff) && (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff));
  assign when_SuperResolutionPart1_l363 = (diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart1_l366 = (diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart1_l371 = ((inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff) && (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff));
  assign when_SuperResolutionPart1_l372 = (diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart1_l375 = (diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart1_l381 = (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart1_l386 = (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign resultStage_pixelStream_ready = (! resultStage_pixelStream_rValid);
  assign resultStage_pixelStream_s2mPipe_valid = (resultStage_pixelStream_valid || resultStage_pixelStream_rValid);
  assign resultStage_pixelStream_s2mPipe_payload = (resultStage_pixelStream_rValid ? resultStage_pixelStream_rData : resultStage_pixelStream_payload);
  always @(*) begin
    resultStage_pixelStream_s2mPipe_ready = resultStage_resultStream_ready;
    if(when_Stream_l368_26) begin
      resultStage_pixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_26 = (! resultStage_resultStream_valid);
  assign resultStage_resultStream_valid = resultStage_pixelStream_s2mPipe_rValid;
  assign resultStage_resultStream_payload = resultStage_pixelStream_s2mPipe_rData;
  assign CICC1851_resultStage_mainOnePixelStream_ready_2 = (CICC1851_resultStage_mainOnePixelStream_ready && CICC1851_resultStage_mainOnePixelStream_ready_1);
  assign CICC1851_resultStage_mainOnePixelStream_ready = (((((resultStage_resultStream_valid && resultStage_mainOnePixelStream_valid) && resultStage_counterOnePixelStream_valid) && resultStage_mainTwoPixelStream_valid) && resultStage_counterTwoPixelStream_valid) && resultStage_controlPipe_valid);
  assign resultStage_resultStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_mainOnePixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_counterOnePixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_mainTwoPixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_counterTwoPixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_controlPipe_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign when_Stream_l438 = (((! resultStage_controlPipe_payload_passValid) && (! resultStage_controlPipe_payload_onceValid)) && (! resultStage_controlPipe_payload_twiceCompValid));
  always @(*) begin
    resultsJoin_valid = CICC1851_resultStage_mainOnePixelStream_ready;
    if(when_Stream_l438) begin
      resultsJoin_valid = 1'b0;
    end
  end

  always @(*) begin
    CICC1851_resultStage_mainOnePixelStream_ready_1 = resultsJoin_ready;
    if(when_Stream_l438) begin
      CICC1851_resultStage_mainOnePixelStream_ready_1 = 1'b1;
    end
  end

  assign pixelsStream_valid = resultsJoin_valid;
  assign resultsJoin_ready = pixelsStream_ready;
  assign pixelsStream_payload_pixel = resultStage_resultStream_payload;
  assign pixelsStream_payload_frameStart = resultStage_controlPipe_payload_frameStart;
  assign pixelsStream_payload_rowEnd = resultStage_controlPipe_payload_rowEnd;
  assign pixelsStream_ready = (! pixelsStream_rValid);
  assign pixelsStream_s2mPipe_valid = (pixelsStream_valid || pixelsStream_rValid);
  assign pixelsStream_s2mPipe_payload_pixel = (pixelsStream_rValid ? pixelsStream_rData_pixel : pixelsStream_payload_pixel);
  assign pixelsStream_s2mPipe_payload_frameStart = (pixelsStream_rValid ? pixelsStream_rData_frameStart : pixelsStream_payload_frameStart);
  assign pixelsStream_s2mPipe_payload_rowEnd = (pixelsStream_rValid ? pixelsStream_rData_rowEnd : pixelsStream_payload_rowEnd);
  always @(*) begin
    pixelsStream_s2mPipe_ready = pixelsStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_27) begin
      pixelsStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_27 = (! pixelsStream_s2mPipe_m2sPipe_valid);
  assign pixelsStream_s2mPipe_m2sPipe_valid = pixelsStream_s2mPipe_rValid;
  assign pixelsStream_s2mPipe_m2sPipe_payload_pixel = pixelsStream_s2mPipe_rData_pixel;
  assign pixelsStream_s2mPipe_m2sPipe_payload_frameStart = pixelsStream_s2mPipe_rData_frameStart;
  assign pixelsStream_s2mPipe_m2sPipe_payload_rowEnd = pixelsStream_s2mPipe_rData_rowEnd;
  assign pixelsStream_s2mPipe_m2sPipe_ready = pixelsOut_ready;
  assign pixelsIn_s2mPipe_valid = (pixelsIn_valid || pixelsIn_rValid);
  assign pixelsIn_s2mPipe_payload_pixel = (pixelsIn_rValid ? pixelsIn_rData_pixel : pixelsIn_payload_pixel);
  assign pixelsIn_s2mPipe_payload_frameStart = (pixelsIn_rValid ? pixelsIn_rData_frameStart : pixelsIn_payload_frameStart);
  assign pixelsIn_s2mPipe_payload_rowEnd = (pixelsIn_rValid ? pixelsIn_rData_rowEnd : pixelsIn_payload_rowEnd);
  always @(*) begin
    pixelsIn_s2mPipe_ready = pixelsIn_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_28) begin
      pixelsIn_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_28 = (! pixelsIn_s2mPipe_m2sPipe_valid);
  assign pixelsIn_s2mPipe_m2sPipe_valid = pixelsIn_s2mPipe_rValid;
  assign pixelsIn_s2mPipe_m2sPipe_payload_pixel = pixelsIn_s2mPipe_rData_pixel;
  assign pixelsIn_s2mPipe_m2sPipe_payload_frameStart = pixelsIn_s2mPipe_rData_frameStart;
  assign pixelsIn_s2mPipe_m2sPipe_payload_rowEnd = pixelsIn_s2mPipe_rData_rowEnd;
  assign passPixels_valid = (pixelsIn_s2mPipe_m2sPipe_valid && bufferEnable);
  assign pixelsIn_s2mPipe_m2sPipe_ready = (passPixels_ready && bufferEnable);
  assign passPixels_payload_pixel = pixelsIn_s2mPipe_m2sPipe_payload_pixel;
  assign passPixels_payload_frameStart = pixelsIn_s2mPipe_m2sPipe_payload_frameStart;
  assign passPixels_payload_rowEnd = pixelsIn_s2mPipe_m2sPipe_payload_rowEnd;
  assign passPixels_ready = 1'b1;
  assign passPixels_fire = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart1_l421 = ((bufferWAddr_value == CICC1851_when_SuperResolutionPart1_l421) && passPixels_fire);
  assign passPixels_fire_1 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart1_l422 = (((bufferRowCount_value == CICC1851_when_SuperResolutionPart1_l422) && bufferReachRowEnd) && passPixels_fire_1);
  assign passPixels_fire_2 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart1_l425 = (passPixels_payload_rowEnd && passPixels_fire_2);
  assign passPixels_fire_3 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart1_l438 = (passPixels_payload_rowEnd && passPixels_fire_3);
  assign passPixels_fire_4 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart1_l439 = (((bufferRowCount_value != 10'h0) && passPixels_payload_rowEnd) && passPixels_fire_4);
  assign when_SuperResolutionPart1_l442 = (bufferReachFinalRow && bufferReachRowEnd);
  assign controlStream_fire = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l447 = (((CICC1851_when_SuperResolutionPart1_l447 == 11'h001) && controlStream_payload_rowEnd) && controlStream_fire);
  assign when_SuperResolutionPart1_l449 = 1'b1;
  assign passPixels_fire_5 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart1_l453 = (passPixels_payload_frameStart && passPixels_fire_5);
  assign passPixels_fire_6 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_7 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_8 = (passPixels_valid && passPixels_ready);
  assign controlStateMachine_wantExit = 1'b0;
  always @(*) begin
    controlStateMachine_wantStart = 1'b0;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_6_HOLD : begin
      end
      controlStateMachine_enumDef_6_PASS : begin
      end
      controlStateMachine_enumDef_6_ONCE : begin
      end
      controlStateMachine_enumDef_6_TWICE : begin
      end
      default : begin
        controlStateMachine_wantStart = 1'b1;
      end
    endcase
  end

  assign controlStateMachine_wantKill = 1'b0;
  always @(*) begin
    controlStateMachine_stateNext = controlStateMachine_stateReg;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_6_HOLD : begin
        if(when_SuperResolutionPart1_l482) begin
          if(passPixels_fire_9) begin
            if(when_SuperResolutionPart1_l484) begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_6_PASS;
            end else begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_6_ONCE;
            end
          end
        end else begin
          if(passPixels_fire_10) begin
            if(when_SuperResolutionPart1_l489) begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_6_ONCE;
            end else begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_6_TWICE;
            end
          end
        end
      end
      controlStateMachine_enumDef_6_PASS : begin
        if(controlStream_fire_1) begin
          if(when_SuperResolutionPart1_l498) begin
            controlStateMachine_stateNext = controlStateMachine_enumDef_6_ONCE;
          end else begin
            if(when_SuperResolutionPart1_l500) begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_6_HOLD;
            end else begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_6_ONCE;
            end
          end
        end
      end
      controlStateMachine_enumDef_6_ONCE : begin
        if(when_SuperResolutionPart1_l537) begin
          if(controlStream_fire_7) begin
            if(outReachRowEnd) begin
              if(bufferReuse) begin
                controlStateMachine_stateNext = controlStateMachine_enumDef_6_ONCE;
              end else begin
                if(when_SuperResolutionPart1_l542) begin
                  controlStateMachine_stateNext = controlStateMachine_enumDef_6_HOLD;
                end else begin
                  controlStateMachine_stateNext = controlStateMachine_enumDef_6_ONCE;
                end
              end
            end else begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_6_PASS;
            end
          end
        end else begin
          if(controlStream_fire_8) begin
            if(bufferReuse) begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_6_TWICE;
            end else begin
              if(when_SuperResolutionPart1_l563) begin
                controlStateMachine_stateNext = controlStateMachine_enumDef_6_HOLD;
              end else begin
                controlStateMachine_stateNext = controlStateMachine_enumDef_6_TWICE;
              end
            end
          end
        end
      end
      controlStateMachine_enumDef_6_TWICE : begin
        if(controlStream_fire_13) begin
          if(outReachRowEnd) begin
            if(bufferReuse) begin
              if(outReachFinalRow) begin
                controlStateMachine_stateNext = controlStateMachine_enumDef_6_HOLD;
              end else begin
                controlStateMachine_stateNext = controlStateMachine_enumDef_6_PASS;
              end
            end else begin
              if(when_SuperResolutionPart1_l612) begin
                controlStateMachine_stateNext = controlStateMachine_enumDef_6_HOLD;
              end else begin
                controlStateMachine_stateNext = controlStateMachine_enumDef_6_PASS;
              end
            end
          end else begin
            controlStateMachine_stateNext = controlStateMachine_enumDef_6_ONCE;
          end
        end
      end
      default : begin
      end
    endcase
    if(controlStateMachine_wantStart) begin
      controlStateMachine_stateNext = controlStateMachine_enumDef_6_HOLD;
    end
    if(controlStateMachine_wantKill) begin
      controlStateMachine_stateNext = controlStateMachine_enumDef_6_BOOT;
    end
  end

  assign when_SuperResolutionPart1_l482 = (CICC1851_when_SuperResolutionPart1_l482 == 11'h0);
  assign passPixels_fire_9 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart1_l484 = (CICC1851_when_SuperResolutionPart1_l484 == 11'h0);
  assign passPixels_fire_10 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart1_l489 = (CICC1851_when_SuperResolutionPart1_l489 == 11'h0);
  assign controlStream_fire_1 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l498 = ((CICC1851_when_SuperResolutionPart1_l498 < CICC1851_when_SuperResolutionPart1_l498_1) || bufferReuse);
  assign passPixels_fire_11 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart1_l500 = ((CICC1851_when_SuperResolutionPart1_l500 == CICC1851_when_SuperResolutionPart1_l500_1) && (! passPixels_fire_11));
  assign controlStream_fire_2 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l507 = (frameStart && controlStream_fire_2);
  assign controlStream_fire_3 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l510 = (controlStream_fire_3 && (CICC1851_when_SuperResolutionPart1_l510 == CICC1851_when_SuperResolutionPart1_l510_1));
  assign controlStream_fire_4 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l511 = ((outReachRowEnd && (CICC1851_when_SuperResolutionPart1_l511 == CICC1851_when_SuperResolutionPart1_l511_1)) && controlStream_fire_4);
  assign controlStream_fire_5 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l513 = (controlStream_fire_5 && outReachRowEnd);
  assign controlStream_fire_6 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l537 = (CICC1851_when_SuperResolutionPart1_l537 == 11'h0);
  assign controlStream_fire_7 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l542 = ((bufferWAddr_value == 10'h0) && (CICC1851_when_SuperResolutionPart1_l542 == CICC1851_when_SuperResolutionPart1_l542_2));
  assign controlStream_fire_8 = (controlStream_valid && controlStream_ready);
  assign passPixels_fire_12 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart1_l563 = ((CICC1851_when_SuperResolutionPart1_l563 == CICC1851_when_SuperResolutionPart1_l563_1) && (! passPixels_fire_12));
  assign controlStream_fire_9 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l578 = (controlStream_fire_9 && (CICC1851_when_SuperResolutionPart1_l578 == CICC1851_when_SuperResolutionPart1_l578_1));
  assign controlStream_fire_10 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l579 = ((outReachRowEnd && (CICC1851_when_SuperResolutionPart1_l579 == CICC1851_when_SuperResolutionPart1_l579_1)) && controlStream_fire_10);
  assign controlStream_fire_11 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l581 = (controlStream_fire_11 && outReachRowEnd);
  assign controlStream_fire_12 = (controlStream_valid && controlStream_ready);
  assign controlStream_fire_13 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l612 = (bufferWAddr_value == 10'h0);
  assign controlStream_fire_14 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l664 = (controlStream_fire_14 && (CICC1851_when_SuperResolutionPart1_l664 == CICC1851_when_SuperResolutionPart1_l664_1));
  assign controlStream_fire_15 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l665 = ((outReachRowEnd && (CICC1851_when_SuperResolutionPart1_l665 == CICC1851_when_SuperResolutionPart1_l665_1)) && controlStream_fire_15);
  assign controlStream_fire_16 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l667 = (controlStream_fire_16 && outReachRowEnd);
  assign controlStream_fire_17 = (controlStream_valid && controlStream_ready);
  always @(posedge clk or negedge resetn) begin
    if(!resetn) begin
      inpDone <= 1'b0;
      readDone <= 1'b0;
      startRead <= 1'b0;
      slaveStart <= 1'b0;
      frameStart <= 1'b0;
      inpThreshold <= 8'h80;
      bmpWidth <= 10'h3c0;
      bmpHeight <= 10'h21c;
      holdBuffer <= 1'b0;
      writeDone <= 1'b0;
      bufferRowCount_value <= 10'h0;
      bufferEnable <= 1'b0;
      bufferSwitch <= 1'b0;
      nextRowBuffer <= 1'b1;
      bufferReuse <= 1'b0;
      bufferWAddr_value <= 10'h0;
      outPixelAddr_value <= 11'h0;
      outRowCount_value <= 11'h0;
      outReachRowEnd <= 1'b0;
      outReachFinalRow <= 1'b0;
      bufferReachRowEnd <= 1'b0;
      bufferReachFinalRow <= 1'b0;
      mainAddrOneStream_rValid <= 1'b0;
      mainAddrOneStream_s2mPipe_rValid <= 1'b0;
      CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_mainOnePixelStream_valid <= 1'b0;
      counterAddrOneStream_rValid <= 1'b0;
      counterAddrOneStream_s2mPipe_rValid <= 1'b0;
      CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_counterOnePixelStream_valid <= 1'b0;
      mainAddrTwoStream_rValid <= 1'b0;
      mainAddrTwoStream_s2mPipe_rValid <= 1'b0;
      CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_mainTwoPixelStream_valid <= 1'b0;
      counterAddrTwoStream_rValid <= 1'b0;
      counterAddrTwoStream_s2mPipe_rValid <= 1'b0;
      CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_counterTwoPixelStream_valid <= 1'b0;
      controlStream_rValid <= 1'b0;
      controlStream_s2mPipe_rValid <= 1'b0;
      controlStream_s2mPipe_m2sPipe_rValid <= 1'b0;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rValid <= 1'b0;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rValid <= 1'b0;
      readStage_mainOnePixelStream_rValid <= 1'b0;
      readStage_mainOnePixelStream_s2mPipe_rValid <= 1'b0;
      readStage_counterOnePixelStream_rValid <= 1'b0;
      readStage_counterOnePixelStream_s2mPipe_rValid <= 1'b0;
      readStage_mainTwoPixelStream_rValid <= 1'b0;
      readStage_mainTwoPixelStream_s2mPipe_rValid <= 1'b0;
      readStage_counterTwoPixelStream_rValid <= 1'b0;
      readStage_counterTwoPixelStream_s2mPipe_rValid <= 1'b0;
      readStage_controlPipe_translated_rValid <= 1'b0;
      readStage_controlPipe_translated_s2mPipe_rValid <= 1'b0;
      compareStage_mainOnePixelStream_rValid <= 1'b0;
      compareStage_mainOnePixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_counterOnePixelStream_rValid <= 1'b0;
      compareStage_counterOnePixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_mainTwoPixelStream_rValid <= 1'b0;
      compareStage_mainTwoPixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_counterTwoPixelStream_rValid <= 1'b0;
      compareStage_counterTwoPixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_controlPipe_translated_rValid <= 1'b0;
      compareStage_controlPipe_translated_s2mPipe_rValid <= 1'b0;
      diffStage_mainOnePixelStream_rValid <= 1'b0;
      diffStage_mainOnePixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_counterOnePixelStream_rValid <= 1'b0;
      diffStage_counterOnePixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_mainTwoPixelStream_rValid <= 1'b0;
      diffStage_mainTwoPixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_counterTwoPixelStream_rValid <= 1'b0;
      diffStage_counterTwoPixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_controlPipe_fork_io_outputs_0_rValid <= 1'b0;
      diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rValid <= 1'b0;
      resultStage_pixelStream_rValid <= 1'b0;
      resultStage_pixelStream_s2mPipe_rValid <= 1'b0;
      pixelsStream_rValid <= 1'b0;
      pixelsStream_s2mPipe_rValid <= 1'b0;
      pixelsIn_rValid <= 1'b0;
      pixelsIn_s2mPipe_rValid <= 1'b0;
      controlStateMachine_stateReg <= controlStateMachine_enumDef_6_BOOT;
    end else begin
      if(when_SuperResolutionPart1_l79) begin
        inpDone <= 1'b1;
      end
      if(when_SuperResolutionPart1_l79_1) begin
        inpDone <= 1'b0;
      end
      if(when_SuperResolutionPart1_l82) begin
        readDone <= 1'b0;
      end
      if(when_SuperResolutionPart1_l85) begin
        startRead <= 1'b1;
      end
      if(when_SuperResolutionPart1_l85_1) begin
        startRead <= 1'b0;
      end
      if(when_SuperResolutionPart1_l88) begin
        slaveStart <= 1'b1;
      end
      if(when_SuperResolutionPart1_l88_1) begin
        slaveStart <= 1'b0;
      end
      inpThreshold <= thresholdIn;
      bmpWidth <= widthIn;
      bmpHeight <= heightIn;
      if(when_SuperResolutionPart1_l103) begin
        holdBuffer <= 1'b0;
      end
      if(when_SuperResolutionPart1_l106) begin
        writeDone <= 1'b0;
      end
      bufferRowCount_value <= bufferRowCount_valueNext;
      if(when_SuperResolutionPart1_l112) begin
        bufferEnable <= 1'b1;
      end
      if(when_SuperResolutionPart1_l112_1) begin
        bufferEnable <= 1'b0;
      end
      if(when_SuperResolutionPart1_l115) begin
        bufferSwitch <= 1'b0;
      end
      if(when_SuperResolutionPart1_l118) begin
        nextRowBuffer <= 1'b1;
      end
      if(inpDone) begin
        bufferReuse <= 1'b0;
      end
      bufferWAddr_value <= bufferWAddr_valueNext;
      outPixelAddr_value <= outPixelAddr_valueNext;
      outRowCount_value <= outRowCount_valueNext;
      if(mainAddrOneStream_valid) begin
        mainAddrOneStream_rValid <= 1'b1;
      end
      if(mainAddrOneStream_s2mPipe_ready) begin
        mainAddrOneStream_rValid <= 1'b0;
      end
      if(mainAddrOneStream_s2mPipe_ready) begin
        mainAddrOneStream_s2mPipe_rValid <= mainAddrOneStream_s2mPipe_valid;
      end
      if(CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(mainAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_2 <= mainAddrOneStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_1) begin
        CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_1) begin
        CICC1851_readStage_mainOnePixelStream_valid <= (CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready || CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_3);
      end
      if(counterAddrOneStream_valid) begin
        counterAddrOneStream_rValid <= 1'b1;
      end
      if(counterAddrOneStream_s2mPipe_ready) begin
        counterAddrOneStream_rValid <= 1'b0;
      end
      if(counterAddrOneStream_s2mPipe_ready) begin
        counterAddrOneStream_s2mPipe_rValid <= counterAddrOneStream_s2mPipe_valid;
      end
      if(CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(counterAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_2 <= counterAddrOneStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_2) begin
        CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_2) begin
        CICC1851_readStage_counterOnePixelStream_valid <= (CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready || CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_3);
      end
      if(mainAddrTwoStream_valid) begin
        mainAddrTwoStream_rValid <= 1'b1;
      end
      if(mainAddrTwoStream_s2mPipe_ready) begin
        mainAddrTwoStream_rValid <= 1'b0;
      end
      if(mainAddrTwoStream_s2mPipe_ready) begin
        mainAddrTwoStream_s2mPipe_rValid <= mainAddrTwoStream_s2mPipe_valid;
      end
      if(CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(mainAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= mainAddrTwoStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_3) begin
        CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_3) begin
        CICC1851_readStage_mainTwoPixelStream_valid <= (CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready || CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_3);
      end
      if(counterAddrTwoStream_valid) begin
        counterAddrTwoStream_rValid <= 1'b1;
      end
      if(counterAddrTwoStream_s2mPipe_ready) begin
        counterAddrTwoStream_rValid <= 1'b0;
      end
      if(counterAddrTwoStream_s2mPipe_ready) begin
        counterAddrTwoStream_s2mPipe_rValid <= counterAddrTwoStream_s2mPipe_valid;
      end
      if(CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(counterAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= counterAddrTwoStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_4) begin
        CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_4) begin
        CICC1851_readStage_counterTwoPixelStream_valid <= (CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready || CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_3);
      end
      if(controlStream_valid) begin
        controlStream_rValid <= 1'b1;
      end
      if(controlStream_s2mPipe_ready) begin
        controlStream_rValid <= 1'b0;
      end
      if(controlStream_s2mPipe_ready) begin
        controlStream_s2mPipe_rValid <= controlStream_s2mPipe_valid;
      end
      if(controlStream_s2mPipe_m2sPipe_ready) begin
        controlStream_s2mPipe_m2sPipe_rValid <= controlStream_s2mPipe_m2sPipe_valid;
      end
      if(controlStream_s2mPipe_m2sPipe_m2sPipe_valid) begin
        controlStream_s2mPipe_m2sPipe_m2sPipe_rValid <= 1'b1;
      end
      if(controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready) begin
        controlStream_s2mPipe_m2sPipe_m2sPipe_rValid <= 1'b0;
      end
      if(controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready) begin
        controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_valid;
      end
      if(readStage_mainOnePixelStream_valid) begin
        readStage_mainOnePixelStream_rValid <= 1'b1;
      end
      if(readStage_mainOnePixelStream_s2mPipe_ready) begin
        readStage_mainOnePixelStream_rValid <= 1'b0;
      end
      if(readStage_mainOnePixelStream_s2mPipe_ready) begin
        readStage_mainOnePixelStream_s2mPipe_rValid <= readStage_mainOnePixelStream_s2mPipe_valid;
      end
      if(readStage_counterOnePixelStream_valid) begin
        readStage_counterOnePixelStream_rValid <= 1'b1;
      end
      if(readStage_counterOnePixelStream_s2mPipe_ready) begin
        readStage_counterOnePixelStream_rValid <= 1'b0;
      end
      if(readStage_counterOnePixelStream_s2mPipe_ready) begin
        readStage_counterOnePixelStream_s2mPipe_rValid <= readStage_counterOnePixelStream_s2mPipe_valid;
      end
      if(readStage_mainTwoPixelStream_valid) begin
        readStage_mainTwoPixelStream_rValid <= 1'b1;
      end
      if(readStage_mainTwoPixelStream_s2mPipe_ready) begin
        readStage_mainTwoPixelStream_rValid <= 1'b0;
      end
      if(readStage_mainTwoPixelStream_s2mPipe_ready) begin
        readStage_mainTwoPixelStream_s2mPipe_rValid <= readStage_mainTwoPixelStream_s2mPipe_valid;
      end
      if(readStage_counterTwoPixelStream_valid) begin
        readStage_counterTwoPixelStream_rValid <= 1'b1;
      end
      if(readStage_counterTwoPixelStream_s2mPipe_ready) begin
        readStage_counterTwoPixelStream_rValid <= 1'b0;
      end
      if(readStage_counterTwoPixelStream_s2mPipe_ready) begin
        readStage_counterTwoPixelStream_s2mPipe_rValid <= readStage_counterTwoPixelStream_s2mPipe_valid;
      end
      if(readStage_controlPipe_translated_valid) begin
        readStage_controlPipe_translated_rValid <= 1'b1;
      end
      if(readStage_controlPipe_translated_s2mPipe_ready) begin
        readStage_controlPipe_translated_rValid <= 1'b0;
      end
      if(readStage_controlPipe_translated_s2mPipe_ready) begin
        readStage_controlPipe_translated_s2mPipe_rValid <= readStage_controlPipe_translated_s2mPipe_valid;
      end
      if(compareStage_mainOnePixelStream_valid) begin
        compareStage_mainOnePixelStream_rValid <= 1'b1;
      end
      if(compareStage_mainOnePixelStream_s2mPipe_ready) begin
        compareStage_mainOnePixelStream_rValid <= 1'b0;
      end
      if(compareStage_mainOnePixelStream_s2mPipe_ready) begin
        compareStage_mainOnePixelStream_s2mPipe_rValid <= compareStage_mainOnePixelStream_s2mPipe_valid;
      end
      if(compareStage_counterOnePixelStream_valid) begin
        compareStage_counterOnePixelStream_rValid <= 1'b1;
      end
      if(compareStage_counterOnePixelStream_s2mPipe_ready) begin
        compareStage_counterOnePixelStream_rValid <= 1'b0;
      end
      if(compareStage_counterOnePixelStream_s2mPipe_ready) begin
        compareStage_counterOnePixelStream_s2mPipe_rValid <= compareStage_counterOnePixelStream_s2mPipe_valid;
      end
      if(compareStage_mainTwoPixelStream_valid) begin
        compareStage_mainTwoPixelStream_rValid <= 1'b1;
      end
      if(compareStage_mainTwoPixelStream_s2mPipe_ready) begin
        compareStage_mainTwoPixelStream_rValid <= 1'b0;
      end
      if(compareStage_mainTwoPixelStream_s2mPipe_ready) begin
        compareStage_mainTwoPixelStream_s2mPipe_rValid <= compareStage_mainTwoPixelStream_s2mPipe_valid;
      end
      if(compareStage_counterTwoPixelStream_valid) begin
        compareStage_counterTwoPixelStream_rValid <= 1'b1;
      end
      if(compareStage_counterTwoPixelStream_s2mPipe_ready) begin
        compareStage_counterTwoPixelStream_rValid <= 1'b0;
      end
      if(compareStage_counterTwoPixelStream_s2mPipe_ready) begin
        compareStage_counterTwoPixelStream_s2mPipe_rValid <= compareStage_counterTwoPixelStream_s2mPipe_valid;
      end
      if(compareStage_controlPipe_translated_valid) begin
        compareStage_controlPipe_translated_rValid <= 1'b1;
      end
      if(compareStage_controlPipe_translated_s2mPipe_ready) begin
        compareStage_controlPipe_translated_rValid <= 1'b0;
      end
      if(compareStage_controlPipe_translated_s2mPipe_ready) begin
        compareStage_controlPipe_translated_s2mPipe_rValid <= compareStage_controlPipe_translated_s2mPipe_valid;
      end
      if(diffStage_mainOnePixelStream_valid) begin
        diffStage_mainOnePixelStream_rValid <= 1'b1;
      end
      if(diffStage_mainOnePixelStream_s2mPipe_ready) begin
        diffStage_mainOnePixelStream_rValid <= 1'b0;
      end
      if(diffStage_mainOnePixelStream_s2mPipe_ready) begin
        diffStage_mainOnePixelStream_s2mPipe_rValid <= diffStage_mainOnePixelStream_s2mPipe_valid;
      end
      if(diffStage_counterOnePixelStream_valid) begin
        diffStage_counterOnePixelStream_rValid <= 1'b1;
      end
      if(diffStage_counterOnePixelStream_s2mPipe_ready) begin
        diffStage_counterOnePixelStream_rValid <= 1'b0;
      end
      if(diffStage_counterOnePixelStream_s2mPipe_ready) begin
        diffStage_counterOnePixelStream_s2mPipe_rValid <= diffStage_counterOnePixelStream_s2mPipe_valid;
      end
      if(diffStage_mainTwoPixelStream_valid) begin
        diffStage_mainTwoPixelStream_rValid <= 1'b1;
      end
      if(diffStage_mainTwoPixelStream_s2mPipe_ready) begin
        diffStage_mainTwoPixelStream_rValid <= 1'b0;
      end
      if(diffStage_mainTwoPixelStream_s2mPipe_ready) begin
        diffStage_mainTwoPixelStream_s2mPipe_rValid <= diffStage_mainTwoPixelStream_s2mPipe_valid;
      end
      if(diffStage_counterTwoPixelStream_valid) begin
        diffStage_counterTwoPixelStream_rValid <= 1'b1;
      end
      if(diffStage_counterTwoPixelStream_s2mPipe_ready) begin
        diffStage_counterTwoPixelStream_rValid <= 1'b0;
      end
      if(diffStage_counterTwoPixelStream_s2mPipe_ready) begin
        diffStage_counterTwoPixelStream_s2mPipe_rValid <= diffStage_counterTwoPixelStream_s2mPipe_valid;
      end
      if(diffStage_controlPipe_fork_io_outputs_0_valid) begin
        diffStage_controlPipe_fork_io_outputs_0_rValid <= 1'b1;
      end
      if(diffStage_controlPipe_fork_io_outputs_0_s2mPipe_ready) begin
        diffStage_controlPipe_fork_io_outputs_0_rValid <= 1'b0;
      end
      if(diffStage_controlPipe_fork_io_outputs_0_s2mPipe_ready) begin
        diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rValid <= diffStage_controlPipe_fork_io_outputs_0_s2mPipe_valid;
      end
      if(resultStage_pixelStream_valid) begin
        resultStage_pixelStream_rValid <= 1'b1;
      end
      if(resultStage_pixelStream_s2mPipe_ready) begin
        resultStage_pixelStream_rValid <= 1'b0;
      end
      if(resultStage_pixelStream_s2mPipe_ready) begin
        resultStage_pixelStream_s2mPipe_rValid <= resultStage_pixelStream_s2mPipe_valid;
      end
      if(pixelsStream_valid) begin
        pixelsStream_rValid <= 1'b1;
      end
      if(pixelsStream_s2mPipe_ready) begin
        pixelsStream_rValid <= 1'b0;
      end
      if(pixelsStream_s2mPipe_ready) begin
        pixelsStream_s2mPipe_rValid <= pixelsStream_s2mPipe_valid;
      end
      if(pixelsIn_valid) begin
        pixelsIn_rValid <= 1'b1;
      end
      if(pixelsIn_s2mPipe_ready) begin
        pixelsIn_rValid <= 1'b0;
      end
      if(pixelsIn_s2mPipe_ready) begin
        pixelsIn_s2mPipe_rValid <= pixelsIn_s2mPipe_valid;
      end
      if(when_SuperResolutionPart1_l421) begin
        bufferReachRowEnd <= 1'b1;
      end
      if(when_SuperResolutionPart1_l422) begin
        bufferReachFinalRow <= 1'b1;
      end
      if(when_SuperResolutionPart1_l425) begin
        if(bufferReachFinalRow) begin
          bufferReuse <= 1'b1;
          bufferReachRowEnd <= 1'b0;
          bufferReachFinalRow <= 1'b0;
        end else begin
          bufferReachRowEnd <= 1'b0;
        end
      end
      if(when_SuperResolutionPart1_l438) begin
        bufferSwitch <= (! bufferSwitch);
      end
      if(when_SuperResolutionPart1_l439) begin
        holdBuffer <= 1'b1;
        bufferEnable <= 1'b0;
        if(when_SuperResolutionPart1_l442) begin
          writeDone <= 1'b1;
          bufferEnable <= 1'b0;
        end
      end
      if(when_SuperResolutionPart1_l447) begin
        holdBuffer <= 1'b0;
        if(when_SuperResolutionPart1_l449) begin
          nextRowBuffer <= (! nextRowBuffer);
        end
      end
      if(when_SuperResolutionPart1_l453) begin
        frameStart <= 1'b1;
      end
      if(inpDone) begin
        inpDone <= 1'b0;
      end
      controlStateMachine_stateReg <= controlStateMachine_stateNext;
      case(controlStateMachine_stateReg)
        controlStateMachine_enumDef_6_HOLD : begin
        end
        controlStateMachine_enumDef_6_PASS : begin
          if(when_SuperResolutionPart1_l507) begin
            frameStart <= 1'b0;
          end
          if(when_SuperResolutionPart1_l510) begin
            outReachRowEnd <= 1'b1;
          end
          if(when_SuperResolutionPart1_l511) begin
            outReachFinalRow <= 1'b1;
          end
          if(when_SuperResolutionPart1_l513) begin
            if(outReachFinalRow) begin
              startRead <= 1'b0;
              readDone <= 1'b1;
              outReachRowEnd <= 1'b0;
              outReachFinalRow <= 1'b0;
            end else begin
              outReachRowEnd <= 1'b0;
            end
          end
          if(controlStream_fire_6) begin
            if(outReachRowEnd) begin
              outReachRowEnd <= 1'b0;
            end
          end
        end
        controlStateMachine_enumDef_6_ONCE : begin
          if(when_SuperResolutionPart1_l578) begin
            outReachRowEnd <= 1'b1;
          end
          if(when_SuperResolutionPart1_l579) begin
            outReachFinalRow <= 1'b1;
          end
          if(when_SuperResolutionPart1_l581) begin
            if(outReachFinalRow) begin
              startRead <= 1'b0;
              readDone <= 1'b1;
              outReachRowEnd <= 1'b0;
              outReachFinalRow <= 1'b0;
            end else begin
              outReachRowEnd <= 1'b0;
            end
          end
          if(controlStream_fire_12) begin
            if(outReachRowEnd) begin
              outReachRowEnd <= 1'b0;
            end
          end
        end
        controlStateMachine_enumDef_6_TWICE : begin
          if(when_SuperResolutionPart1_l664) begin
            outReachRowEnd <= 1'b1;
          end
          if(when_SuperResolutionPart1_l665) begin
            outReachFinalRow <= 1'b1;
          end
          if(when_SuperResolutionPart1_l667) begin
            if(outReachFinalRow) begin
              startRead <= 1'b0;
              readDone <= 1'b1;
              outReachRowEnd <= 1'b0;
              outReachFinalRow <= 1'b0;
            end else begin
              outReachRowEnd <= 1'b0;
            end
          end
          if(controlStream_fire_17) begin
            if(outReachRowEnd) begin
              outReachRowEnd <= 1'b0;
            end
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(posedge clk) begin
    startIn_regNext <= startIn;
    if(mainAddrOneStream_ready) begin
      mainAddrOneStream_rData <= mainAddrOneStream_payload;
    end
    if(mainAddrOneStream_s2mPipe_ready) begin
      mainAddrOneStream_s2mPipe_rData <= mainAddrOneStream_s2mPipe_payload;
    end
    if(CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_mainOnePixelStream_payload_1 <= CICC1851_readStage_mainOnePixelStream_payload;
    end
    if(CICC1851_1) begin
      CICC1851_readStage_mainOnePixelStream_payload_2 <= (CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_mainOnePixelStream_payload_1 : CICC1851_readStage_mainOnePixelStream_payload);
    end
    if(counterAddrOneStream_ready) begin
      counterAddrOneStream_rData <= counterAddrOneStream_payload;
    end
    if(counterAddrOneStream_s2mPipe_ready) begin
      counterAddrOneStream_s2mPipe_rData <= counterAddrOneStream_s2mPipe_payload;
    end
    if(CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_counterOnePixelStream_payload_1 <= CICC1851_readStage_counterOnePixelStream_payload;
    end
    if(CICC1851_2) begin
      CICC1851_readStage_counterOnePixelStream_payload_2 <= (CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_counterOnePixelStream_payload_1 : CICC1851_readStage_counterOnePixelStream_payload);
    end
    if(mainAddrTwoStream_ready) begin
      mainAddrTwoStream_rData <= mainAddrTwoStream_payload;
    end
    if(mainAddrTwoStream_s2mPipe_ready) begin
      mainAddrTwoStream_s2mPipe_rData <= mainAddrTwoStream_s2mPipe_payload;
    end
    if(CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_mainTwoPixelStream_payload_1 <= CICC1851_readStage_mainTwoPixelStream_payload;
    end
    if(CICC1851_3) begin
      CICC1851_readStage_mainTwoPixelStream_payload_2 <= (CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_mainTwoPixelStream_payload_1 : CICC1851_readStage_mainTwoPixelStream_payload);
    end
    if(counterAddrTwoStream_ready) begin
      counterAddrTwoStream_rData <= counterAddrTwoStream_payload;
    end
    if(counterAddrTwoStream_s2mPipe_ready) begin
      counterAddrTwoStream_s2mPipe_rData <= counterAddrTwoStream_s2mPipe_payload;
    end
    if(CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_counterTwoPixelStream_payload_1 <= CICC1851_readStage_counterTwoPixelStream_payload;
    end
    if(CICC1851_4) begin
      CICC1851_readStage_counterTwoPixelStream_payload_2 <= (CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_counterTwoPixelStream_payload_1 : CICC1851_readStage_counterTwoPixelStream_payload);
    end
    if(controlStream_ready) begin
      controlStream_rData_frameStart <= controlStream_payload_frameStart;
      controlStream_rData_rowEnd <= controlStream_payload_rowEnd;
      controlStream_rData_passMode <= controlStream_payload_passMode;
      controlStream_rData_passValid <= controlStream_payload_passValid;
      controlStream_rData_onceMode <= controlStream_payload_onceMode;
      controlStream_rData_onceValid <= controlStream_payload_onceValid;
      controlStream_rData_mainCompare <= controlStream_payload_mainCompare;
      controlStream_rData_counterCompare <= controlStream_payload_counterCompare;
      controlStream_rData_mainDiff <= controlStream_payload_mainDiff;
      controlStream_rData_counterDiff <= controlStream_payload_counterDiff;
      controlStream_rData_twiceCompValid <= controlStream_payload_twiceCompValid;
      controlStream_rData_twiceMode <= controlStream_payload_twiceMode;
    end
    if(controlStream_s2mPipe_ready) begin
      controlStream_s2mPipe_rData_frameStart <= controlStream_s2mPipe_payload_frameStart;
      controlStream_s2mPipe_rData_rowEnd <= controlStream_s2mPipe_payload_rowEnd;
      controlStream_s2mPipe_rData_passMode <= controlStream_s2mPipe_payload_passMode;
      controlStream_s2mPipe_rData_passValid <= controlStream_s2mPipe_payload_passValid;
      controlStream_s2mPipe_rData_onceMode <= controlStream_s2mPipe_payload_onceMode;
      controlStream_s2mPipe_rData_onceValid <= controlStream_s2mPipe_payload_onceValid;
      controlStream_s2mPipe_rData_mainCompare <= controlStream_s2mPipe_payload_mainCompare;
      controlStream_s2mPipe_rData_counterCompare <= controlStream_s2mPipe_payload_counterCompare;
      controlStream_s2mPipe_rData_mainDiff <= controlStream_s2mPipe_payload_mainDiff;
      controlStream_s2mPipe_rData_counterDiff <= controlStream_s2mPipe_payload_counterDiff;
      controlStream_s2mPipe_rData_twiceCompValid <= controlStream_s2mPipe_payload_twiceCompValid;
      controlStream_s2mPipe_rData_twiceMode <= controlStream_s2mPipe_payload_twiceMode;
    end
    if(controlStream_s2mPipe_m2sPipe_ready) begin
      controlStream_s2mPipe_m2sPipe_rData_frameStart <= controlStream_s2mPipe_m2sPipe_payload_frameStart;
      controlStream_s2mPipe_m2sPipe_rData_rowEnd <= controlStream_s2mPipe_m2sPipe_payload_rowEnd;
      controlStream_s2mPipe_m2sPipe_rData_passMode <= controlStream_s2mPipe_m2sPipe_payload_passMode;
      controlStream_s2mPipe_m2sPipe_rData_passValid <= controlStream_s2mPipe_m2sPipe_payload_passValid;
      controlStream_s2mPipe_m2sPipe_rData_onceMode <= controlStream_s2mPipe_m2sPipe_payload_onceMode;
      controlStream_s2mPipe_m2sPipe_rData_onceValid <= controlStream_s2mPipe_m2sPipe_payload_onceValid;
      controlStream_s2mPipe_m2sPipe_rData_mainCompare <= controlStream_s2mPipe_m2sPipe_payload_mainCompare;
      controlStream_s2mPipe_m2sPipe_rData_counterCompare <= controlStream_s2mPipe_m2sPipe_payload_counterCompare;
      controlStream_s2mPipe_m2sPipe_rData_mainDiff <= controlStream_s2mPipe_m2sPipe_payload_mainDiff;
      controlStream_s2mPipe_m2sPipe_rData_counterDiff <= controlStream_s2mPipe_m2sPipe_payload_counterDiff;
      controlStream_s2mPipe_m2sPipe_rData_twiceCompValid <= controlStream_s2mPipe_m2sPipe_payload_twiceCompValid;
      controlStream_s2mPipe_m2sPipe_rData_twiceMode <= controlStream_s2mPipe_m2sPipe_payload_twiceMode;
    end
    if(controlStream_s2mPipe_m2sPipe_m2sPipe_ready) begin
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_frameStart <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_frameStart;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_rowEnd <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_rowEnd;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_passMode <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passMode;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_passValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_onceMode <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceMode;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_onceValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_twiceCompValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceCompValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_twiceMode <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceMode;
    end
    if(controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready) begin
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_frameStart <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_frameStart;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_rowEnd <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_rowEnd;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_passMode <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_passMode;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_passValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_passValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_onceMode <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_onceMode;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_onceValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_onceValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_twiceCompValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_twiceCompValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_twiceMode <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_twiceMode;
    end
    if(readStage_mainOnePixelStream_ready) begin
      readStage_mainOnePixelStream_rData <= readStage_mainOnePixelStream_payload;
    end
    if(readStage_mainOnePixelStream_s2mPipe_ready) begin
      readStage_mainOnePixelStream_s2mPipe_rData <= readStage_mainOnePixelStream_s2mPipe_payload;
    end
    if(readStage_counterOnePixelStream_ready) begin
      readStage_counterOnePixelStream_rData <= readStage_counterOnePixelStream_payload;
    end
    if(readStage_counterOnePixelStream_s2mPipe_ready) begin
      readStage_counterOnePixelStream_s2mPipe_rData <= readStage_counterOnePixelStream_s2mPipe_payload;
    end
    if(readStage_mainTwoPixelStream_ready) begin
      readStage_mainTwoPixelStream_rData <= readStage_mainTwoPixelStream_payload;
    end
    if(readStage_mainTwoPixelStream_s2mPipe_ready) begin
      readStage_mainTwoPixelStream_s2mPipe_rData <= readStage_mainTwoPixelStream_s2mPipe_payload;
    end
    if(readStage_counterTwoPixelStream_ready) begin
      readStage_counterTwoPixelStream_rData <= readStage_counterTwoPixelStream_payload;
    end
    if(readStage_counterTwoPixelStream_s2mPipe_ready) begin
      readStage_counterTwoPixelStream_s2mPipe_rData <= readStage_counterTwoPixelStream_s2mPipe_payload;
    end
    if(readStage_controlPipe_translated_ready) begin
      readStage_controlPipe_translated_rData_frameStart <= readStage_controlPipe_translated_payload_frameStart;
      readStage_controlPipe_translated_rData_rowEnd <= readStage_controlPipe_translated_payload_rowEnd;
      readStage_controlPipe_translated_rData_passMode <= readStage_controlPipe_translated_payload_passMode;
      readStage_controlPipe_translated_rData_passValid <= readStage_controlPipe_translated_payload_passValid;
      readStage_controlPipe_translated_rData_onceMode <= readStage_controlPipe_translated_payload_onceMode;
      readStage_controlPipe_translated_rData_onceValid <= readStage_controlPipe_translated_payload_onceValid;
      readStage_controlPipe_translated_rData_mainCompare <= readStage_controlPipe_translated_payload_mainCompare;
      readStage_controlPipe_translated_rData_counterCompare <= readStage_controlPipe_translated_payload_counterCompare;
      readStage_controlPipe_translated_rData_mainDiff <= readStage_controlPipe_translated_payload_mainDiff;
      readStage_controlPipe_translated_rData_counterDiff <= readStage_controlPipe_translated_payload_counterDiff;
      readStage_controlPipe_translated_rData_twiceCompValid <= readStage_controlPipe_translated_payload_twiceCompValid;
      readStage_controlPipe_translated_rData_twiceMode <= readStage_controlPipe_translated_payload_twiceMode;
    end
    if(readStage_controlPipe_translated_s2mPipe_ready) begin
      readStage_controlPipe_translated_s2mPipe_rData_frameStart <= readStage_controlPipe_translated_s2mPipe_payload_frameStart;
      readStage_controlPipe_translated_s2mPipe_rData_rowEnd <= readStage_controlPipe_translated_s2mPipe_payload_rowEnd;
      readStage_controlPipe_translated_s2mPipe_rData_passMode <= readStage_controlPipe_translated_s2mPipe_payload_passMode;
      readStage_controlPipe_translated_s2mPipe_rData_passValid <= readStage_controlPipe_translated_s2mPipe_payload_passValid;
      readStage_controlPipe_translated_s2mPipe_rData_onceMode <= readStage_controlPipe_translated_s2mPipe_payload_onceMode;
      readStage_controlPipe_translated_s2mPipe_rData_onceValid <= readStage_controlPipe_translated_s2mPipe_payload_onceValid;
      readStage_controlPipe_translated_s2mPipe_rData_mainCompare <= readStage_controlPipe_translated_s2mPipe_payload_mainCompare;
      readStage_controlPipe_translated_s2mPipe_rData_counterCompare <= readStage_controlPipe_translated_s2mPipe_payload_counterCompare;
      readStage_controlPipe_translated_s2mPipe_rData_mainDiff <= readStage_controlPipe_translated_s2mPipe_payload_mainDiff;
      readStage_controlPipe_translated_s2mPipe_rData_counterDiff <= readStage_controlPipe_translated_s2mPipe_payload_counterDiff;
      readStage_controlPipe_translated_s2mPipe_rData_twiceCompValid <= readStage_controlPipe_translated_s2mPipe_payload_twiceCompValid;
      readStage_controlPipe_translated_s2mPipe_rData_twiceMode <= readStage_controlPipe_translated_s2mPipe_payload_twiceMode;
    end
    if(compareStage_mainOnePixelStream_ready) begin
      compareStage_mainOnePixelStream_rData <= compareStage_mainOnePixelStream_payload;
    end
    if(compareStage_mainOnePixelStream_s2mPipe_ready) begin
      compareStage_mainOnePixelStream_s2mPipe_rData <= compareStage_mainOnePixelStream_s2mPipe_payload;
    end
    if(compareStage_counterOnePixelStream_ready) begin
      compareStage_counterOnePixelStream_rData <= compareStage_counterOnePixelStream_payload;
    end
    if(compareStage_counterOnePixelStream_s2mPipe_ready) begin
      compareStage_counterOnePixelStream_s2mPipe_rData <= compareStage_counterOnePixelStream_s2mPipe_payload;
    end
    if(compareStage_mainTwoPixelStream_ready) begin
      compareStage_mainTwoPixelStream_rData <= compareStage_mainTwoPixelStream_payload;
    end
    if(compareStage_mainTwoPixelStream_s2mPipe_ready) begin
      compareStage_mainTwoPixelStream_s2mPipe_rData <= compareStage_mainTwoPixelStream_s2mPipe_payload;
    end
    if(compareStage_counterTwoPixelStream_ready) begin
      compareStage_counterTwoPixelStream_rData <= compareStage_counterTwoPixelStream_payload;
    end
    if(compareStage_counterTwoPixelStream_s2mPipe_ready) begin
      compareStage_counterTwoPixelStream_s2mPipe_rData <= compareStage_counterTwoPixelStream_s2mPipe_payload;
    end
    if(compareStage_controlPipe_translated_ready) begin
      compareStage_controlPipe_translated_rData_frameStart <= compareStage_controlPipe_translated_payload_frameStart;
      compareStage_controlPipe_translated_rData_rowEnd <= compareStage_controlPipe_translated_payload_rowEnd;
      compareStage_controlPipe_translated_rData_passMode <= compareStage_controlPipe_translated_payload_passMode;
      compareStage_controlPipe_translated_rData_passValid <= compareStage_controlPipe_translated_payload_passValid;
      compareStage_controlPipe_translated_rData_onceMode <= compareStage_controlPipe_translated_payload_onceMode;
      compareStage_controlPipe_translated_rData_onceValid <= compareStage_controlPipe_translated_payload_onceValid;
      compareStage_controlPipe_translated_rData_mainCompare <= compareStage_controlPipe_translated_payload_mainCompare;
      compareStage_controlPipe_translated_rData_counterCompare <= compareStage_controlPipe_translated_payload_counterCompare;
      compareStage_controlPipe_translated_rData_mainDiff <= compareStage_controlPipe_translated_payload_mainDiff;
      compareStage_controlPipe_translated_rData_counterDiff <= compareStage_controlPipe_translated_payload_counterDiff;
      compareStage_controlPipe_translated_rData_twiceCompValid <= compareStage_controlPipe_translated_payload_twiceCompValid;
      compareStage_controlPipe_translated_rData_twiceMode <= compareStage_controlPipe_translated_payload_twiceMode;
    end
    if(compareStage_controlPipe_translated_s2mPipe_ready) begin
      compareStage_controlPipe_translated_s2mPipe_rData_frameStart <= compareStage_controlPipe_translated_s2mPipe_payload_frameStart;
      compareStage_controlPipe_translated_s2mPipe_rData_rowEnd <= compareStage_controlPipe_translated_s2mPipe_payload_rowEnd;
      compareStage_controlPipe_translated_s2mPipe_rData_passMode <= compareStage_controlPipe_translated_s2mPipe_payload_passMode;
      compareStage_controlPipe_translated_s2mPipe_rData_passValid <= compareStage_controlPipe_translated_s2mPipe_payload_passValid;
      compareStage_controlPipe_translated_s2mPipe_rData_onceMode <= compareStage_controlPipe_translated_s2mPipe_payload_onceMode;
      compareStage_controlPipe_translated_s2mPipe_rData_onceValid <= compareStage_controlPipe_translated_s2mPipe_payload_onceValid;
      compareStage_controlPipe_translated_s2mPipe_rData_mainCompare <= compareStage_controlPipe_translated_s2mPipe_payload_mainCompare;
      compareStage_controlPipe_translated_s2mPipe_rData_counterCompare <= compareStage_controlPipe_translated_s2mPipe_payload_counterCompare;
      compareStage_controlPipe_translated_s2mPipe_rData_mainDiff <= compareStage_controlPipe_translated_s2mPipe_payload_mainDiff;
      compareStage_controlPipe_translated_s2mPipe_rData_counterDiff <= compareStage_controlPipe_translated_s2mPipe_payload_counterDiff;
      compareStage_controlPipe_translated_s2mPipe_rData_twiceCompValid <= compareStage_controlPipe_translated_s2mPipe_payload_twiceCompValid;
      compareStage_controlPipe_translated_s2mPipe_rData_twiceMode <= compareStage_controlPipe_translated_s2mPipe_payload_twiceMode;
    end
    if(diffStage_mainOnePixelStream_ready) begin
      diffStage_mainOnePixelStream_rData <= diffStage_mainOnePixelStream_payload;
    end
    if(diffStage_mainOnePixelStream_s2mPipe_ready) begin
      diffStage_mainOnePixelStream_s2mPipe_rData <= diffStage_mainOnePixelStream_s2mPipe_payload;
    end
    if(diffStage_counterOnePixelStream_ready) begin
      diffStage_counterOnePixelStream_rData <= diffStage_counterOnePixelStream_payload;
    end
    if(diffStage_counterOnePixelStream_s2mPipe_ready) begin
      diffStage_counterOnePixelStream_s2mPipe_rData <= diffStage_counterOnePixelStream_s2mPipe_payload;
    end
    if(diffStage_mainTwoPixelStream_ready) begin
      diffStage_mainTwoPixelStream_rData <= diffStage_mainTwoPixelStream_payload;
    end
    if(diffStage_mainTwoPixelStream_s2mPipe_ready) begin
      diffStage_mainTwoPixelStream_s2mPipe_rData <= diffStage_mainTwoPixelStream_s2mPipe_payload;
    end
    if(diffStage_counterTwoPixelStream_ready) begin
      diffStage_counterTwoPixelStream_rData <= diffStage_counterTwoPixelStream_payload;
    end
    if(diffStage_counterTwoPixelStream_s2mPipe_ready) begin
      diffStage_counterTwoPixelStream_s2mPipe_rData <= diffStage_counterTwoPixelStream_s2mPipe_payload;
    end
    if(diffStage_controlPipe_fork_io_outputs_0_ready) begin
      diffStage_controlPipe_fork_io_outputs_0_rData_frameStart <= diffStage_controlPipe_fork_io_outputs_0_payload_frameStart;
      diffStage_controlPipe_fork_io_outputs_0_rData_rowEnd <= diffStage_controlPipe_fork_io_outputs_0_payload_rowEnd;
      diffStage_controlPipe_fork_io_outputs_0_rData_passMode <= diffStage_controlPipe_fork_io_outputs_0_payload_passMode;
      diffStage_controlPipe_fork_io_outputs_0_rData_passValid <= diffStage_controlPipe_fork_io_outputs_0_payload_passValid;
      diffStage_controlPipe_fork_io_outputs_0_rData_onceMode <= diffStage_controlPipe_fork_io_outputs_0_payload_onceMode;
      diffStage_controlPipe_fork_io_outputs_0_rData_onceValid <= diffStage_controlPipe_fork_io_outputs_0_payload_onceValid;
      diffStage_controlPipe_fork_io_outputs_0_rData_mainCompare <= diffStage_controlPipe_fork_io_outputs_0_payload_mainCompare;
      diffStage_controlPipe_fork_io_outputs_0_rData_counterCompare <= diffStage_controlPipe_fork_io_outputs_0_payload_counterCompare;
      diffStage_controlPipe_fork_io_outputs_0_rData_mainDiff <= diffStage_controlPipe_fork_io_outputs_0_payload_mainDiff;
      diffStage_controlPipe_fork_io_outputs_0_rData_counterDiff <= diffStage_controlPipe_fork_io_outputs_0_payload_counterDiff;
      diffStage_controlPipe_fork_io_outputs_0_rData_twiceCompValid <= diffStage_controlPipe_fork_io_outputs_0_payload_twiceCompValid;
      diffStage_controlPipe_fork_io_outputs_0_rData_twiceMode <= diffStage_controlPipe_fork_io_outputs_0_payload_twiceMode;
    end
    if(diffStage_controlPipe_fork_io_outputs_0_s2mPipe_ready) begin
      diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_frameStart <= diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_frameStart;
      diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_rowEnd <= diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_rowEnd;
      diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_passMode <= diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_passMode;
      diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_passValid <= diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_passValid;
      diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_onceMode <= diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_onceMode;
      diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_onceValid <= diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_onceValid;
      diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_mainCompare <= diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_mainCompare;
      diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_counterCompare <= diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_counterCompare;
      diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_mainDiff <= diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_mainDiff;
      diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_counterDiff <= diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_counterDiff;
      diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_twiceCompValid <= diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_twiceCompValid;
      diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_twiceMode <= diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_twiceMode;
    end
    if(resultStage_pixelStream_ready) begin
      resultStage_pixelStream_rData <= resultStage_pixelStream_payload;
    end
    if(resultStage_pixelStream_s2mPipe_ready) begin
      resultStage_pixelStream_s2mPipe_rData <= resultStage_pixelStream_s2mPipe_payload;
    end
    if(pixelsStream_ready) begin
      pixelsStream_rData_pixel <= pixelsStream_payload_pixel;
      pixelsStream_rData_frameStart <= pixelsStream_payload_frameStart;
      pixelsStream_rData_rowEnd <= pixelsStream_payload_rowEnd;
    end
    if(pixelsStream_s2mPipe_ready) begin
      pixelsStream_s2mPipe_rData_pixel <= pixelsStream_s2mPipe_payload_pixel;
      pixelsStream_s2mPipe_rData_frameStart <= pixelsStream_s2mPipe_payload_frameStart;
      pixelsStream_s2mPipe_rData_rowEnd <= pixelsStream_s2mPipe_payload_rowEnd;
    end
    if(pixelsIn_ready) begin
      pixelsIn_rData_pixel <= pixelsIn_payload_pixel;
      pixelsIn_rData_frameStart <= pixelsIn_payload_frameStart;
      pixelsIn_rData_rowEnd <= pixelsIn_payload_rowEnd;
    end
    if(pixelsIn_s2mPipe_ready) begin
      pixelsIn_s2mPipe_rData_pixel <= pixelsIn_s2mPipe_payload_pixel;
      pixelsIn_s2mPipe_rData_frameStart <= pixelsIn_s2mPipe_payload_frameStart;
      pixelsIn_s2mPipe_rData_rowEnd <= pixelsIn_s2mPipe_payload_rowEnd;
    end
  end


endmodule

module SuperResolutionPart3_1 (
  input               pixelsIn_valid,
  output reg          pixelsIn_ready,
  input      [7:0]    pixelsIn_payload_pixel,
  input               pixelsIn_payload_frameStart,
  input               pixelsIn_payload_rowEnd,
  input               pixelsIn_payload_inpValid,
  input               startIn,
  output reg          pixelsOut_valid,
  input               pixelsOut_ready,
  output reg [7:0]    pixelsOut_payload_pixel,
  output reg          pixelsOut_payload_frameStart,
  output reg          pixelsOut_payload_rowEnd,
  output reg          inpThreeDoneOut,
  input      [7:0]    thresholdIn,
  input      [9:0]    widthIn,
  input      [9:0]    heightIn,
  input               clk,
  input               resetn
);
  localparam controlStateMachine_enumDef_5_BOOT = 2'd0;
  localparam controlStateMachine_enumDef_5_HOLD = 2'd1;
  localparam controlStateMachine_enumDef_5_PASS = 2'd2;
  localparam controlStateMachine_enumDef_5_EXTRA = 2'd3;

  reg        [7:0]    CICC1851_lineBufferOne_port1;
  reg        [7:0]    CICC1851_lineBufferOne_port2;
  reg        [7:0]    CICC1851_lineBufferTwo_port1;
  reg        [7:0]    CICC1851_lineBufferTwo_port2;
  reg        [7:0]    CICC1851_lineBufferThree_port1;
  reg        [7:0]    CICC1851_lineBufferThree_port2;
  reg        [0:0]    CICC1851_validBufferOne_port1;
  reg        [0:0]    CICC1851_validBufferOne_port2;
  reg        [0:0]    CICC1851_validBufferTwo_port1;
  reg        [0:0]    CICC1851_validBufferTwo_port2;
  reg        [0:0]    CICC1851_validBufferThree_port1;
  reg        [0:0]    CICC1851_validBufferThree_port2;
  wire                diffStage_controlPipe_fork_io_input_ready;
  wire                diffStage_controlPipe_fork_io_outputs_0_valid;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_frameStart;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_rowEnd;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_pipeValid;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_firstRow;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_lastRow;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_finalResult;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_mainCompare;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_counterCompare;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_horizontalCompare;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_verticalCompare;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_payload_mainDiff;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_payload_counterDiff;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_payload_horizontalDiff;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_payload_verticalDiff;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_isHorizontalMin;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_payload_minDiff;
  wire       [1:0]    diffStage_controlPipe_fork_io_outputs_0_payload_currentPosition;
  wire       [1:0]    diffStage_controlPipe_fork_io_outputs_0_payload_nextPosition;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_horizontalDirectionValid;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_verticalDirectionValid;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_mainDirectionValid;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_counterDirectionValid;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_inValidMinDiff;
  wire                diffStage_controlPipe_fork_io_outputs_1_valid;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_frameStart;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_rowEnd;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_pipeValid;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_firstRow;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_lastRow;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_finalResult;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_mainCompare;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_counterCompare;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_horizontalCompare;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_verticalCompare;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_1_payload_horizontalDiff;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_1_payload_verticalDiff;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_isHorizontalMin;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_1_payload_minDiff;
  wire       [1:0]    diffStage_controlPipe_fork_io_outputs_1_payload_currentPosition;
  wire       [1:0]    diffStage_controlPipe_fork_io_outputs_1_payload_nextPosition;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_horizontalDirectionValid;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_verticalDirectionValid;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_mainDirectionValid;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_counterDirectionValid;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_inValidMinDiff;
  wire       [11:0]   CICC1851_bufferRowCount_valueNext;
  wire       [0:0]    CICC1851_bufferRowCount_valueNext_1;
  wire       [11:0]   CICC1851_bufferWAddr_valueNext;
  wire       [0:0]    CICC1851_bufferWAddr_valueNext_1;
  wire       [11:0]   CICC1851_outPixelAddr_valueNext;
  wire       [0:0]    CICC1851_outPixelAddr_valueNext_1;
  wire       [11:0]   CICC1851_outRowCount_valueNext;
  wire       [0:0]    CICC1851_outRowCount_valueNext_1;
  wire       [11:0]   CICC1851_alreadySendRow_valueNext;
  wire       [0:0]    CICC1851_alreadySendRow_valueNext_1;
  wire       [11:0]   CICC1851_alreadySendCountInRow_valueNext;
  wire       [0:0]    CICC1851_alreadySendCountInRow_valueNext_1;
  wire       [0:0]    CICC1851_nextRowBuffer;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l226;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l226_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l226_2;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l227;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l227_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l227_2;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l270;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l270_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l270_2;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l271;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l271_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l271_2;
  wire       [7:0]    CICC1851_lineBufferOne_port;
  wire                CICC1851_lineBufferOne_port_1;
  wire       [7:0]    CICC1851_lineBufferTwo_port;
  wire                CICC1851_lineBufferTwo_port_1;
  wire       [7:0]    CICC1851_lineBufferThree_port;
  wire                CICC1851_lineBufferThree_port_1;
  wire       [0:0]    CICC1851_validBufferOne_port;
  wire                CICC1851_validBufferOne_port_1;
  wire       [0:0]    CICC1851_validBufferTwo_port;
  wire                CICC1851_validBufferTwo_port_1;
  wire       [0:0]    CICC1851_validBufferThree_port;
  wire                CICC1851_validBufferThree_port_1;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_1;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_2;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_3;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_4;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_5;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_6;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_7;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_8;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_9;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_10;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_11;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_12;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_13;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_14;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_15;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_16;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_17;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_18;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_19;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_20;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_21;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_22;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_23;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_24;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_25;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_26;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_27;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_28;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_29;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_30;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_31;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_32;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_33;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_34;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_35;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_36;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_37;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_38;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_39;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_40;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_41;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_42;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_43;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_44;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_45;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_46;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_47;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_48;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_49;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_50;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_51;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_52;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_53;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_54;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_55;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_56;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_57;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_58;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_59;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_60;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_61;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_62;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_63;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_64;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_65;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_66;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_67;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_68;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_69;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_70;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_71;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_72;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_73;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_74;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_75;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_76;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_77;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_78;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_79;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_80;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_81;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_82;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_83;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_84;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_85;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_86;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_87;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_88;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_89;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_90;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_91;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_92;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_93;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_94;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_95;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_96;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_97;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_98;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_99;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_100;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_101;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_102;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_103;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_104;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_105;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_106;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_107;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_108;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_109;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_110;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_111;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_112;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_113;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_114;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_115;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_116;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_117;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_118;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_119;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_120;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_121;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_122;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_123;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_124;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_125;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_126;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_127;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_128;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_129;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_130;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_131;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_132;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_133;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_134;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_135;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_136;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_137;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_138;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_139;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_140;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_141;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_142;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_143;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_144;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_145;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_146;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_147;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_148;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_149;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_150;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_151;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_152;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_153;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_154;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_155;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_156;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_157;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_158;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_159;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_160;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_161;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_162;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_163;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_164;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_165;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_166;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_167;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_168;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_169;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_170;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_171;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_172;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_173;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_174;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_175;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_176;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_177;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_178;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_179;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_180;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_181;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_182;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_183;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_184;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_185;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_186;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_187;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_188;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_189;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_190;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_191;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_192;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_193;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_194;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_195;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_196;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_197;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_198;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_199;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_200;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_201;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_202;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_203;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_204;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_205;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_206;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_207;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_208;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_209;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_210;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_211;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_212;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_213;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_214;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_215;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_216;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_217;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_218;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_219;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_220;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_221;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_222;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_223;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_224;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_225;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_226;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_227;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_228;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_229;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_230;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_231;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_232;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_233;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_234;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_235;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_236;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_237;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_238;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_239;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_240;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_241;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_242;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_243;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_244;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_245;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_246;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_247;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_248;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_249;
  wire       [11:0]   CICC1851_when_SuperResolutionPart3_l1202;
  wire       [11:0]   CICC1851_when_SuperResolutionPart3_l1205;
  wire       [11:0]   CICC1851_when_SuperResolutionPart3_l1205_1;
  wire       [11:0]   CICC1851_when_SuperResolutionPart3_l1205_2;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l1223;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l1223_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l1223_2;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l1224;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l1224_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l1224_2;
  reg                 inpThreeDone;
  reg                 startIn_regNext;
  wire                when_SuperResolutionPart3_l72;
  reg                 readDone;
  wire                when_SuperResolutionPart3_l75;
  reg                 startRead;
  wire                when_SuperResolutionPart3_l78;
  wire                when_SuperResolutionPart3_l78_1;
  reg                 frameStart;
  reg        [7:0]    inpThreshold;
  reg        [9:0]    bmpWidth;
  reg        [9:0]    bmpHeight;
  reg                 holdBuffer;
  wire                when_SuperResolutionPart3_l93;
  reg                 writeDone;
  wire                when_SuperResolutionPart3_l96;
  reg                 bufferRowCount_willIncrement;
  reg                 bufferRowCount_willClear;
  reg        [11:0]   bufferRowCount_valueNext;
  reg        [11:0]   bufferRowCount_value;
  wire                bufferRowCount_willOverflowIfInc;
  wire                bufferRowCount_willOverflow;
  reg                 bufferEnable;
  wire                when_SuperResolutionPart3_l102;
  wire                when_SuperResolutionPart3_l102_1;
  reg        [1:0]    bufferSwitch;
  reg        [1:0]    nextRowBuffer;
  reg        [1:0]    currentRowBuffer;
  reg                 bufferReuse;
  reg                 bufferWAddr_willIncrement;
  reg                 bufferWAddr_willClear;
  reg        [11:0]   bufferWAddr_valueNext;
  reg        [11:0]   bufferWAddr_value;
  wire                bufferWAddr_willOverflowIfInc;
  wire                bufferWAddr_willOverflow;
  reg                 outPixelAddr_willIncrement;
  reg                 outPixelAddr_willClear;
  reg        [11:0]   outPixelAddr_valueNext;
  reg        [11:0]   outPixelAddr_value;
  wire                outPixelAddr_willOverflowIfInc;
  wire                outPixelAddr_willOverflow;
  reg                 outRowCount_willIncrement;
  reg                 outRowCount_willClear;
  reg        [11:0]   outRowCount_valueNext;
  reg        [11:0]   outRowCount_value;
  wire                outRowCount_willOverflowIfInc;
  wire                outRowCount_willOverflow;
  reg                 alreadySendRow_willIncrement;
  reg                 alreadySendRow_willClear;
  reg        [11:0]   alreadySendRow_valueNext;
  reg        [11:0]   alreadySendRow_value;
  wire                alreadySendRow_willOverflowIfInc;
  wire                alreadySendRow_willOverflow;
  reg                 alreadySendCountInRow_willIncrement;
  reg                 alreadySendCountInRow_willClear;
  reg        [11:0]   alreadySendCountInRow_valueNext;
  reg        [11:0]   alreadySendCountInRow_value;
  wire                alreadySendCountInRow_willOverflowIfInc;
  wire                alreadySendCountInRow_willOverflow;
  reg                 alreadyReachRowEnd;
  reg                 alreadyReachFinalRow;
  reg                 outReachRowEnd;
  reg                 outReachFinalRow;
  reg                 bufferReachRowEnd;
  reg                 bufferReachFinalRow;
  reg        [7:0]    minDiff;
  reg        [7:0]    candidatePixel;
  reg                 isHorizontalDirection;
  reg                 inValidMinDiff;
  reg                 startIn_regNext_1;
  wire                when_SuperResolutionPart3_l154;
  reg        [11:0]   mainAddrOne;
  reg        [11:0]   counterAddrOne;
  reg        [11:0]   mainAddrTwo;
  reg        [11:0]   counterAddrTwo;
  reg        [11:0]   mainAddrThree;
  reg        [11:0]   counterAddrThree;
  wire                validStream_valid;
  reg                 validStream_ready;
  wire                controlStream_valid;
  wire                controlStream_ready;
  wire                controlStream_payload_frameStart;
  wire                controlStream_payload_rowEnd;
  wire                controlStream_payload_pipeValid;
  wire                controlStream_payload_firstRow;
  wire                controlStream_payload_lastRow;
  wire                controlStream_payload_finalResult;
  wire                controlStream_payload_mainCompare;
  wire                controlStream_payload_counterCompare;
  wire                controlStream_payload_horizontalCompare;
  wire                controlStream_payload_verticalCompare;
  wire       [7:0]    controlStream_payload_mainDiff;
  wire       [7:0]    controlStream_payload_counterDiff;
  wire       [7:0]    controlStream_payload_horizontalDiff;
  wire       [7:0]    controlStream_payload_verticalDiff;
  wire                controlStream_payload_isHorizontalMin;
  wire       [7:0]    controlStream_payload_minDiff;
  wire       [1:0]    controlStream_payload_currentPosition;
  wire       [1:0]    controlStream_payload_nextPosition;
  wire                controlStream_payload_horizontalDirectionValid;
  wire                controlStream_payload_verticalDirectionValid;
  wire                controlStream_payload_mainDirectionValid;
  wire                controlStream_payload_counterDirectionValid;
  wire                controlStream_payload_inValidMinDiff;
  reg                 controls_frameStart;
  reg                 controls_rowEnd;
  reg                 controls_pipeValid;
  reg                 controls_firstRow;
  reg                 controls_lastRow;
  reg                 controls_finalResult;
  wire                controls_mainCompare;
  wire                controls_counterCompare;
  wire                controls_horizontalCompare;
  wire                controls_verticalCompare;
  wire       [7:0]    controls_mainDiff;
  wire       [7:0]    controls_counterDiff;
  wire       [7:0]    controls_horizontalDiff;
  wire       [7:0]    controls_verticalDiff;
  wire                controls_isHorizontalMin;
  wire       [7:0]    controls_minDiff;
  reg        [1:0]    controls_currentPosition;
  reg        [1:0]    controls_nextPosition;
  wire                controls_horizontalDirectionValid;
  wire                controls_verticalDirectionValid;
  wire                controls_mainDirectionValid;
  wire                controls_counterDirectionValid;
  wire                controls_inValidMinDiff;
  wire       [59:0]   CICC1851_controls_frameStart;
  wire                mainPixelAddrOneStream_valid;
  wire                mainPixelAddrOneStream_ready;
  wire       [11:0]   mainPixelAddrOneStream_payload;
  wire                counterPixelAddrOneStream_valid;
  wire                counterPixelAddrOneStream_ready;
  wire       [11:0]   counterPixelAddrOneStream_payload;
  wire                mainPixelAddrTwoStream_valid;
  wire                mainPixelAddrTwoStream_ready;
  wire       [11:0]   mainPixelAddrTwoStream_payload;
  wire                counterPixelAddrTwoStream_valid;
  wire                counterPixelAddrTwoStream_ready;
  wire       [11:0]   counterPixelAddrTwoStream_payload;
  wire                mainPixelAddrThreeStream_valid;
  wire                mainPixelAddrThreeStream_ready;
  wire       [11:0]   mainPixelAddrThreeStream_payload;
  wire                counterPixelAddrThreeStream_valid;
  wire                counterPixelAddrThreeStream_ready;
  wire       [11:0]   counterPixelAddrThreeStream_payload;
  wire                mainValidAddrOneStream_valid;
  wire                mainValidAddrOneStream_ready;
  wire       [11:0]   mainValidAddrOneStream_payload;
  wire                counterValidAddrOneStream_valid;
  wire                counterValidAddrOneStream_ready;
  wire       [11:0]   counterValidAddrOneStream_payload;
  wire                mainValidAddrTwoStream_valid;
  wire                mainValidAddrTwoStream_ready;
  wire       [11:0]   mainValidAddrTwoStream_payload;
  wire                counterValidAddrTwoStream_valid;
  wire                counterValidAddrTwoStream_ready;
  wire       [11:0]   counterValidAddrTwoStream_payload;
  wire                mainValidAddrThreeStream_valid;
  wire                mainValidAddrThreeStream_ready;
  wire       [11:0]   mainValidAddrThreeStream_payload;
  wire                counterValidAddrThreeStream_valid;
  wire                counterValidAddrThreeStream_ready;
  wire       [11:0]   counterValidAddrThreeStream_payload;
  wire                pixelsIn_s2mPipe_valid;
  reg                 pixelsIn_s2mPipe_ready;
  wire       [7:0]    pixelsIn_s2mPipe_payload_pixel;
  wire                pixelsIn_s2mPipe_payload_frameStart;
  wire                pixelsIn_s2mPipe_payload_rowEnd;
  wire                pixelsIn_s2mPipe_payload_inpValid;
  reg                 pixelsIn_rValid;
  reg        [7:0]    pixelsIn_rData_pixel;
  reg                 pixelsIn_rData_frameStart;
  reg                 pixelsIn_rData_rowEnd;
  reg                 pixelsIn_rData_inpValid;
  wire                pixelsIn_s2mPipe_m2sPipe_valid;
  wire                pixelsIn_s2mPipe_m2sPipe_ready;
  wire       [7:0]    pixelsIn_s2mPipe_m2sPipe_payload_pixel;
  wire                pixelsIn_s2mPipe_m2sPipe_payload_frameStart;
  wire                pixelsIn_s2mPipe_m2sPipe_payload_rowEnd;
  wire                pixelsIn_s2mPipe_m2sPipe_payload_inpValid;
  reg                 pixelsIn_s2mPipe_rValid;
  reg        [7:0]    pixelsIn_s2mPipe_rData_pixel;
  reg                 pixelsIn_s2mPipe_rData_frameStart;
  reg                 pixelsIn_s2mPipe_rData_rowEnd;
  reg                 pixelsIn_s2mPipe_rData_inpValid;
  wire                when_Stream_l368;
  wire                passPixels_valid;
  wire                passPixels_ready;
  wire       [7:0]    passPixels_payload_pixel;
  wire                passPixels_payload_frameStart;
  wire                passPixels_payload_rowEnd;
  wire                passPixels_payload_inpValid;
  wire                passPixels_fire;
  wire                when_SuperResolutionPart3_l226;
  wire                passPixels_fire_1;
  wire                when_SuperResolutionPart3_l227;
  wire                passPixels_fire_2;
  wire                when_SuperResolutionPart3_l230;
  wire                passPixels_fire_3;
  wire                when_SuperResolutionPart3_l243;
  wire                when_SuperResolutionPart3_l244;
  wire                passPixels_fire_4;
  wire                when_SuperResolutionPart3_l251;
  wire                when_SuperResolutionPart3_l255;
  wire                passPixels_fire_5;
  wire                when_SuperResolutionPart3_l262;
  wire                pixelsOut_fire;
  wire                when_SuperResolutionPart3_l270;
  wire                pixelsOut_fire_1;
  wire                when_SuperResolutionPart3_l271;
  wire                pixelsOut_fire_2;
  wire                pixelsOut_fire_3;
  wire                when_SuperResolutionPart3_l282;
  wire                passPixels_fire_6;
  wire                passPixels_fire_7;
  wire                passPixels_fire_8;
  wire                passPixels_fire_9;
  wire                passPixels_fire_10;
  wire                passPixels_fire_11;
  wire                passPixels_fire_12;
  wire                mainPixelAddrOneStream_s2mPipe_valid;
  reg                 mainPixelAddrOneStream_s2mPipe_ready;
  wire       [11:0]   mainPixelAddrOneStream_s2mPipe_payload;
  reg                 mainPixelAddrOneStream_rValid;
  reg        [11:0]   mainPixelAddrOneStream_rData;
  wire                mainPixelAddrOneStream_s2mPipe_m2sPipe_valid;
  wire                mainPixelAddrOneStream_s2mPipe_m2sPipe_ready;
  wire       [11:0]   mainPixelAddrOneStream_s2mPipe_m2sPipe_payload;
  reg                 mainPixelAddrOneStream_s2mPipe_rValid;
  reg        [11:0]   mainPixelAddrOneStream_s2mPipe_rData;
  wire                when_Stream_l368_1;
  wire                CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_mainOnePixelStream_payload;
  reg                 CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_1;
  reg                 CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_mainOnePixelStream_payload_1;
  wire                readStage_mainOnePixelStream_valid;
  wire                readStage_mainOnePixelStream_ready;
  wire       [7:0]    readStage_mainOnePixelStream_payload;
  reg                 CICC1851_readStage_mainOnePixelStream_valid;
  reg        [7:0]    CICC1851_readStage_mainOnePixelStream_payload_2;
  wire                when_Stream_l368_2;
  wire                counterPixelAddrOneStream_s2mPipe_valid;
  reg                 counterPixelAddrOneStream_s2mPipe_ready;
  wire       [11:0]   counterPixelAddrOneStream_s2mPipe_payload;
  reg                 counterPixelAddrOneStream_rValid;
  reg        [11:0]   counterPixelAddrOneStream_rData;
  wire                counterPixelAddrOneStream_s2mPipe_m2sPipe_valid;
  wire                counterPixelAddrOneStream_s2mPipe_m2sPipe_ready;
  wire       [11:0]   counterPixelAddrOneStream_s2mPipe_m2sPipe_payload;
  reg                 counterPixelAddrOneStream_s2mPipe_rValid;
  reg        [11:0]   counterPixelAddrOneStream_s2mPipe_rData;
  wire                when_Stream_l368_3;
  wire                CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_counterOnePixelStream_payload;
  reg                 CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_2;
  reg                 CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_counterOnePixelStream_payload_1;
  wire                readStage_counterOnePixelStream_valid;
  wire                readStage_counterOnePixelStream_ready;
  wire       [7:0]    readStage_counterOnePixelStream_payload;
  reg                 CICC1851_readStage_counterOnePixelStream_valid;
  reg        [7:0]    CICC1851_readStage_counterOnePixelStream_payload_2;
  wire                when_Stream_l368_4;
  wire                mainPixelAddrTwoStream_s2mPipe_valid;
  reg                 mainPixelAddrTwoStream_s2mPipe_ready;
  wire       [11:0]   mainPixelAddrTwoStream_s2mPipe_payload;
  reg                 mainPixelAddrTwoStream_rValid;
  reg        [11:0]   mainPixelAddrTwoStream_rData;
  wire                mainPixelAddrTwoStream_s2mPipe_m2sPipe_valid;
  wire                mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire       [11:0]   mainPixelAddrTwoStream_s2mPipe_m2sPipe_payload;
  reg                 mainPixelAddrTwoStream_s2mPipe_rValid;
  reg        [11:0]   mainPixelAddrTwoStream_s2mPipe_rData;
  wire                when_Stream_l368_5;
  wire                CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_mainTwoPixelStream_payload;
  reg                 CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_3;
  reg                 CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_mainTwoPixelStream_payload_1;
  wire                readStage_mainTwoPixelStream_valid;
  wire                readStage_mainTwoPixelStream_ready;
  wire       [7:0]    readStage_mainTwoPixelStream_payload;
  reg                 CICC1851_readStage_mainTwoPixelStream_valid;
  reg        [7:0]    CICC1851_readStage_mainTwoPixelStream_payload_2;
  wire                when_Stream_l368_6;
  wire                counterPixelAddrTwoStream_s2mPipe_valid;
  reg                 counterPixelAddrTwoStream_s2mPipe_ready;
  wire       [11:0]   counterPixelAddrTwoStream_s2mPipe_payload;
  reg                 counterPixelAddrTwoStream_rValid;
  reg        [11:0]   counterPixelAddrTwoStream_rData;
  wire                counterPixelAddrTwoStream_s2mPipe_m2sPipe_valid;
  wire                counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire       [11:0]   counterPixelAddrTwoStream_s2mPipe_m2sPipe_payload;
  reg                 counterPixelAddrTwoStream_s2mPipe_rValid;
  reg        [11:0]   counterPixelAddrTwoStream_s2mPipe_rData;
  wire                when_Stream_l368_7;
  wire                CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_counterTwoPixelStream_payload;
  reg                 CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_4;
  reg                 CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_counterTwoPixelStream_payload_1;
  wire                readStage_counterTwoPixelStream_valid;
  wire                readStage_counterTwoPixelStream_ready;
  wire       [7:0]    readStage_counterTwoPixelStream_payload;
  reg                 CICC1851_readStage_counterTwoPixelStream_valid;
  reg        [7:0]    CICC1851_readStage_counterTwoPixelStream_payload_2;
  wire                when_Stream_l368_8;
  wire                mainPixelAddrThreeStream_s2mPipe_valid;
  reg                 mainPixelAddrThreeStream_s2mPipe_ready;
  wire       [11:0]   mainPixelAddrThreeStream_s2mPipe_payload;
  reg                 mainPixelAddrThreeStream_rValid;
  reg        [11:0]   mainPixelAddrThreeStream_rData;
  wire                mainPixelAddrThreeStream_s2mPipe_m2sPipe_valid;
  wire                mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready;
  wire       [11:0]   mainPixelAddrThreeStream_s2mPipe_m2sPipe_payload;
  reg                 mainPixelAddrThreeStream_s2mPipe_rValid;
  reg        [11:0]   mainPixelAddrThreeStream_s2mPipe_rData;
  wire                when_Stream_l368_9;
  wire                CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_mainThreePixelStream_payload;
  reg                 CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_5;
  reg                 CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_mainThreePixelStream_payload_1;
  wire                readStage_mainThreePixelStream_valid;
  wire                readStage_mainThreePixelStream_ready;
  wire       [7:0]    readStage_mainThreePixelStream_payload;
  reg                 CICC1851_readStage_mainThreePixelStream_valid;
  reg        [7:0]    CICC1851_readStage_mainThreePixelStream_payload_2;
  wire                when_Stream_l368_10;
  wire                counterPixelAddrThreeStream_s2mPipe_valid;
  reg                 counterPixelAddrThreeStream_s2mPipe_ready;
  wire       [11:0]   counterPixelAddrThreeStream_s2mPipe_payload;
  reg                 counterPixelAddrThreeStream_rValid;
  reg        [11:0]   counterPixelAddrThreeStream_rData;
  wire                counterPixelAddrThreeStream_s2mPipe_m2sPipe_valid;
  wire                counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready;
  wire       [11:0]   counterPixelAddrThreeStream_s2mPipe_m2sPipe_payload;
  reg                 counterPixelAddrThreeStream_s2mPipe_rValid;
  reg        [11:0]   counterPixelAddrThreeStream_s2mPipe_rData;
  wire                when_Stream_l368_11;
  wire                CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_counterThreePixelStream_payload;
  reg                 CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_6;
  reg                 CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_counterThreePixelStream_payload_1;
  wire                readStage_counterThreePixelStream_valid;
  wire                readStage_counterThreePixelStream_ready;
  wire       [7:0]    readStage_counterThreePixelStream_payload;
  reg                 CICC1851_readStage_counterThreePixelStream_valid;
  reg        [7:0]    CICC1851_readStage_counterThreePixelStream_payload_2;
  wire                when_Stream_l368_12;
  wire                mainValidAddrOneStream_s2mPipe_valid;
  reg                 mainValidAddrOneStream_s2mPipe_ready;
  wire       [11:0]   mainValidAddrOneStream_s2mPipe_payload;
  reg                 mainValidAddrOneStream_rValid;
  reg        [11:0]   mainValidAddrOneStream_rData;
  wire                mainValidAddrOneStream_s2mPipe_m2sPipe_valid;
  wire                mainValidAddrOneStream_s2mPipe_m2sPipe_ready;
  wire       [11:0]   mainValidAddrOneStream_s2mPipe_m2sPipe_payload;
  reg                 mainValidAddrOneStream_s2mPipe_rValid;
  reg        [11:0]   mainValidAddrOneStream_s2mPipe_rData;
  wire                when_Stream_l368_13;
  wire                CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_1;
  wire                CICC1851_readStage_mainOneValidStream_payload;
  reg                 CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_7;
  reg                 CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_3;
  reg                 CICC1851_readStage_mainOneValidStream_payload_1;
  wire                readStage_mainOneValidStream_valid;
  wire                readStage_mainOneValidStream_ready;
  wire                readStage_mainOneValidStream_payload;
  reg                 CICC1851_readStage_mainOneValidStream_valid;
  reg                 CICC1851_readStage_mainOneValidStream_payload_2;
  wire                when_Stream_l368_14;
  wire                counterValidAddrOneStream_s2mPipe_valid;
  reg                 counterValidAddrOneStream_s2mPipe_ready;
  wire       [11:0]   counterValidAddrOneStream_s2mPipe_payload;
  reg                 counterValidAddrOneStream_rValid;
  reg        [11:0]   counterValidAddrOneStream_rData;
  wire                counterValidAddrOneStream_s2mPipe_m2sPipe_valid;
  wire                counterValidAddrOneStream_s2mPipe_m2sPipe_ready;
  wire       [11:0]   counterValidAddrOneStream_s2mPipe_m2sPipe_payload;
  reg                 counterValidAddrOneStream_s2mPipe_rValid;
  reg        [11:0]   counterValidAddrOneStream_s2mPipe_rData;
  wire                when_Stream_l368_15;
  wire                CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_1;
  wire                CICC1851_readStage_counterOneValidStream_payload;
  reg                 CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_8;
  reg                 CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_3;
  reg                 CICC1851_readStage_counterOneValidStream_payload_1;
  wire                readStage_counterOneValidStream_valid;
  wire                readStage_counterOneValidStream_ready;
  wire                readStage_counterOneValidStream_payload;
  reg                 CICC1851_readStage_counterOneValidStream_valid;
  reg                 CICC1851_readStage_counterOneValidStream_payload_2;
  wire                when_Stream_l368_16;
  wire                mainValidAddrTwoStream_s2mPipe_valid;
  reg                 mainValidAddrTwoStream_s2mPipe_ready;
  wire       [11:0]   mainValidAddrTwoStream_s2mPipe_payload;
  reg                 mainValidAddrTwoStream_rValid;
  reg        [11:0]   mainValidAddrTwoStream_rData;
  wire                mainValidAddrTwoStream_s2mPipe_m2sPipe_valid;
  wire                mainValidAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire       [11:0]   mainValidAddrTwoStream_s2mPipe_m2sPipe_payload;
  reg                 mainValidAddrTwoStream_s2mPipe_rValid;
  reg        [11:0]   mainValidAddrTwoStream_s2mPipe_rData;
  wire                when_Stream_l368_17;
  wire                CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_1;
  wire                CICC1851_readStage_mainTwoValidStream_payload;
  reg                 CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_9;
  reg                 CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_3;
  reg                 CICC1851_readStage_mainTwoValidStream_payload_1;
  wire                readStage_mainTwoValidStream_valid;
  wire                readStage_mainTwoValidStream_ready;
  wire                readStage_mainTwoValidStream_payload;
  reg                 CICC1851_readStage_mainTwoValidStream_valid;
  reg                 CICC1851_readStage_mainTwoValidStream_payload_2;
  wire                when_Stream_l368_18;
  wire                counterValidAddrTwoStream_s2mPipe_valid;
  reg                 counterValidAddrTwoStream_s2mPipe_ready;
  wire       [11:0]   counterValidAddrTwoStream_s2mPipe_payload;
  reg                 counterValidAddrTwoStream_rValid;
  reg        [11:0]   counterValidAddrTwoStream_rData;
  wire                counterValidAddrTwoStream_s2mPipe_m2sPipe_valid;
  wire                counterValidAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire       [11:0]   counterValidAddrTwoStream_s2mPipe_m2sPipe_payload;
  reg                 counterValidAddrTwoStream_s2mPipe_rValid;
  reg        [11:0]   counterValidAddrTwoStream_s2mPipe_rData;
  wire                when_Stream_l368_19;
  wire                CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_1;
  wire                CICC1851_readStage_counterTwoValidStream_payload;
  reg                 CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_10;
  reg                 CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_3;
  reg                 CICC1851_readStage_counterTwoValidStream_payload_1;
  wire                readStage_counterTwoValidStream_valid;
  wire                readStage_counterTwoValidStream_ready;
  wire                readStage_counterTwoValidStream_payload;
  reg                 CICC1851_readStage_counterTwoValidStream_valid;
  reg                 CICC1851_readStage_counterTwoValidStream_payload_2;
  wire                when_Stream_l368_20;
  wire                mainValidAddrThreeStream_s2mPipe_valid;
  reg                 mainValidAddrThreeStream_s2mPipe_ready;
  wire       [11:0]   mainValidAddrThreeStream_s2mPipe_payload;
  reg                 mainValidAddrThreeStream_rValid;
  reg        [11:0]   mainValidAddrThreeStream_rData;
  wire                mainValidAddrThreeStream_s2mPipe_m2sPipe_valid;
  wire                mainValidAddrThreeStream_s2mPipe_m2sPipe_ready;
  wire       [11:0]   mainValidAddrThreeStream_s2mPipe_m2sPipe_payload;
  reg                 mainValidAddrThreeStream_s2mPipe_rValid;
  reg        [11:0]   mainValidAddrThreeStream_s2mPipe_rData;
  wire                when_Stream_l368_21;
  wire                CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_1;
  wire                CICC1851_readStage_mainThreeValidStream_payload;
  reg                 CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_11;
  reg                 CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_3;
  reg                 CICC1851_readStage_mainThreeValidStream_payload_1;
  wire                readStage_mainThreeValidStream_valid;
  wire                readStage_mainThreeValidStream_ready;
  wire                readStage_mainThreeValidStream_payload;
  reg                 CICC1851_readStage_mainThreeValidStream_valid;
  reg                 CICC1851_readStage_mainThreeValidStream_payload_2;
  wire                when_Stream_l368_22;
  wire                counterValidAddrThreeStream_s2mPipe_valid;
  reg                 counterValidAddrThreeStream_s2mPipe_ready;
  wire       [11:0]   counterValidAddrThreeStream_s2mPipe_payload;
  reg                 counterValidAddrThreeStream_rValid;
  reg        [11:0]   counterValidAddrThreeStream_rData;
  wire                counterValidAddrThreeStream_s2mPipe_m2sPipe_valid;
  wire                counterValidAddrThreeStream_s2mPipe_m2sPipe_ready;
  wire       [11:0]   counterValidAddrThreeStream_s2mPipe_m2sPipe_payload;
  reg                 counterValidAddrThreeStream_s2mPipe_rValid;
  reg        [11:0]   counterValidAddrThreeStream_s2mPipe_rData;
  wire                when_Stream_l368_23;
  wire                CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_1;
  wire                CICC1851_readStage_counterThreeValidStream_payload;
  reg                 CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_12;
  reg                 CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_3;
  reg                 CICC1851_readStage_counterThreeValidStream_payload_1;
  wire                readStage_counterThreeValidStream_valid;
  wire                readStage_counterThreeValidStream_ready;
  wire                readStage_counterThreeValidStream_payload;
  reg                 CICC1851_readStage_counterThreeValidStream_valid;
  reg                 CICC1851_readStage_counterThreeValidStream_payload_2;
  wire                when_Stream_l368_24;
  wire                controlStream_s2mPipe_valid;
  reg                 controlStream_s2mPipe_ready;
  wire                controlStream_s2mPipe_payload_frameStart;
  wire                controlStream_s2mPipe_payload_rowEnd;
  wire                controlStream_s2mPipe_payload_pipeValid;
  wire                controlStream_s2mPipe_payload_firstRow;
  wire                controlStream_s2mPipe_payload_lastRow;
  wire                controlStream_s2mPipe_payload_finalResult;
  wire                controlStream_s2mPipe_payload_mainCompare;
  wire                controlStream_s2mPipe_payload_counterCompare;
  wire                controlStream_s2mPipe_payload_horizontalCompare;
  wire                controlStream_s2mPipe_payload_verticalCompare;
  wire       [7:0]    controlStream_s2mPipe_payload_mainDiff;
  wire       [7:0]    controlStream_s2mPipe_payload_counterDiff;
  wire       [7:0]    controlStream_s2mPipe_payload_horizontalDiff;
  wire       [7:0]    controlStream_s2mPipe_payload_verticalDiff;
  wire                controlStream_s2mPipe_payload_isHorizontalMin;
  wire       [7:0]    controlStream_s2mPipe_payload_minDiff;
  wire       [1:0]    controlStream_s2mPipe_payload_currentPosition;
  wire       [1:0]    controlStream_s2mPipe_payload_nextPosition;
  wire                controlStream_s2mPipe_payload_horizontalDirectionValid;
  wire                controlStream_s2mPipe_payload_verticalDirectionValid;
  wire                controlStream_s2mPipe_payload_mainDirectionValid;
  wire                controlStream_s2mPipe_payload_counterDirectionValid;
  wire                controlStream_s2mPipe_payload_inValidMinDiff;
  reg                 controlStream_rValid;
  reg                 controlStream_rData_frameStart;
  reg                 controlStream_rData_rowEnd;
  reg                 controlStream_rData_pipeValid;
  reg                 controlStream_rData_firstRow;
  reg                 controlStream_rData_lastRow;
  reg                 controlStream_rData_finalResult;
  reg                 controlStream_rData_mainCompare;
  reg                 controlStream_rData_counterCompare;
  reg                 controlStream_rData_horizontalCompare;
  reg                 controlStream_rData_verticalCompare;
  reg        [7:0]    controlStream_rData_mainDiff;
  reg        [7:0]    controlStream_rData_counterDiff;
  reg        [7:0]    controlStream_rData_horizontalDiff;
  reg        [7:0]    controlStream_rData_verticalDiff;
  reg                 controlStream_rData_isHorizontalMin;
  reg        [7:0]    controlStream_rData_minDiff;
  reg        [1:0]    controlStream_rData_currentPosition;
  reg        [1:0]    controlStream_rData_nextPosition;
  reg                 controlStream_rData_horizontalDirectionValid;
  reg                 controlStream_rData_verticalDirectionValid;
  reg                 controlStream_rData_mainDirectionValid;
  reg                 controlStream_rData_counterDirectionValid;
  reg                 controlStream_rData_inValidMinDiff;
  wire                controlStream_s2mPipe_m2sPipe_valid;
  reg                 controlStream_s2mPipe_m2sPipe_ready;
  wire                controlStream_s2mPipe_m2sPipe_payload_frameStart;
  wire                controlStream_s2mPipe_m2sPipe_payload_rowEnd;
  wire                controlStream_s2mPipe_m2sPipe_payload_pipeValid;
  wire                controlStream_s2mPipe_m2sPipe_payload_firstRow;
  wire                controlStream_s2mPipe_m2sPipe_payload_lastRow;
  wire                controlStream_s2mPipe_m2sPipe_payload_finalResult;
  wire                controlStream_s2mPipe_m2sPipe_payload_mainCompare;
  wire                controlStream_s2mPipe_m2sPipe_payload_counterCompare;
  wire                controlStream_s2mPipe_m2sPipe_payload_horizontalCompare;
  wire                controlStream_s2mPipe_m2sPipe_payload_verticalCompare;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_payload_mainDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_payload_counterDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_payload_horizontalDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_payload_verticalDiff;
  wire                controlStream_s2mPipe_m2sPipe_payload_isHorizontalMin;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_payload_minDiff;
  wire       [1:0]    controlStream_s2mPipe_m2sPipe_payload_currentPosition;
  wire       [1:0]    controlStream_s2mPipe_m2sPipe_payload_nextPosition;
  wire                controlStream_s2mPipe_m2sPipe_payload_horizontalDirectionValid;
  wire                controlStream_s2mPipe_m2sPipe_payload_verticalDirectionValid;
  wire                controlStream_s2mPipe_m2sPipe_payload_mainDirectionValid;
  wire                controlStream_s2mPipe_m2sPipe_payload_counterDirectionValid;
  wire                controlStream_s2mPipe_m2sPipe_payload_inValidMinDiff;
  reg                 controlStream_s2mPipe_rValid;
  reg                 controlStream_s2mPipe_rData_frameStart;
  reg                 controlStream_s2mPipe_rData_rowEnd;
  reg                 controlStream_s2mPipe_rData_pipeValid;
  reg                 controlStream_s2mPipe_rData_firstRow;
  reg                 controlStream_s2mPipe_rData_lastRow;
  reg                 controlStream_s2mPipe_rData_finalResult;
  reg                 controlStream_s2mPipe_rData_mainCompare;
  reg                 controlStream_s2mPipe_rData_counterCompare;
  reg                 controlStream_s2mPipe_rData_horizontalCompare;
  reg                 controlStream_s2mPipe_rData_verticalCompare;
  reg        [7:0]    controlStream_s2mPipe_rData_mainDiff;
  reg        [7:0]    controlStream_s2mPipe_rData_counterDiff;
  reg        [7:0]    controlStream_s2mPipe_rData_horizontalDiff;
  reg        [7:0]    controlStream_s2mPipe_rData_verticalDiff;
  reg                 controlStream_s2mPipe_rData_isHorizontalMin;
  reg        [7:0]    controlStream_s2mPipe_rData_minDiff;
  reg        [1:0]    controlStream_s2mPipe_rData_currentPosition;
  reg        [1:0]    controlStream_s2mPipe_rData_nextPosition;
  reg                 controlStream_s2mPipe_rData_horizontalDirectionValid;
  reg                 controlStream_s2mPipe_rData_verticalDirectionValid;
  reg                 controlStream_s2mPipe_rData_mainDirectionValid;
  reg                 controlStream_s2mPipe_rData_counterDirectionValid;
  reg                 controlStream_s2mPipe_rData_inValidMinDiff;
  wire                when_Stream_l368_25;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_valid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_ready;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_frameStart;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_rowEnd;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_pipeValid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_firstRow;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_lastRow;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_finalResult;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainCompare;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterCompare;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_horizontalCompare;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_verticalCompare;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_horizontalDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_verticalDiff;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_isHorizontalMin;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_minDiff;
  wire       [1:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_currentPosition;
  wire       [1:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_nextPosition;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_horizontalDirectionValid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_verticalDirectionValid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDirectionValid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDirectionValid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_inValidMinDiff;
  reg                 controlStream_s2mPipe_m2sPipe_rValid;
  reg                 controlStream_s2mPipe_m2sPipe_rData_frameStart;
  reg                 controlStream_s2mPipe_m2sPipe_rData_rowEnd;
  reg                 controlStream_s2mPipe_m2sPipe_rData_pipeValid;
  reg                 controlStream_s2mPipe_m2sPipe_rData_firstRow;
  reg                 controlStream_s2mPipe_m2sPipe_rData_lastRow;
  reg                 controlStream_s2mPipe_m2sPipe_rData_finalResult;
  reg                 controlStream_s2mPipe_m2sPipe_rData_mainCompare;
  reg                 controlStream_s2mPipe_m2sPipe_rData_counterCompare;
  reg                 controlStream_s2mPipe_m2sPipe_rData_horizontalCompare;
  reg                 controlStream_s2mPipe_m2sPipe_rData_verticalCompare;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_rData_mainDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_rData_counterDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_rData_horizontalDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_rData_verticalDiff;
  reg                 controlStream_s2mPipe_m2sPipe_rData_isHorizontalMin;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_rData_minDiff;
  reg        [1:0]    controlStream_s2mPipe_m2sPipe_rData_currentPosition;
  reg        [1:0]    controlStream_s2mPipe_m2sPipe_rData_nextPosition;
  reg                 controlStream_s2mPipe_m2sPipe_rData_horizontalDirectionValid;
  reg                 controlStream_s2mPipe_m2sPipe_rData_verticalDirectionValid;
  reg                 controlStream_s2mPipe_m2sPipe_rData_mainDirectionValid;
  reg                 controlStream_s2mPipe_m2sPipe_rData_counterDirectionValid;
  reg                 controlStream_s2mPipe_m2sPipe_rData_inValidMinDiff;
  wire                when_Stream_l368_26;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_valid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_frameStart;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_rowEnd;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_pipeValid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_firstRow;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_lastRow;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_finalResult;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainCompare;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterCompare;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_horizontalCompare;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_verticalCompare;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_horizontalDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_verticalDiff;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_isHorizontalMin;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_minDiff;
  wire       [1:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_currentPosition;
  wire       [1:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_nextPosition;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_horizontalDirectionValid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_verticalDirectionValid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainDirectionValid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterDirectionValid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_inValidMinDiff;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_frameStart;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_rowEnd;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_pipeValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_firstRow;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_lastRow;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_finalResult;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainCompare;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterCompare;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_horizontalCompare;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_verticalCompare;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_horizontalDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_verticalDiff;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_isHorizontalMin;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_minDiff;
  reg        [1:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_currentPosition;
  reg        [1:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_nextPosition;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_horizontalDirectionValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_verticalDirectionValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainDirectionValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterDirectionValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_inValidMinDiff;
  wire                readStage_controlPipe_valid;
  wire                readStage_controlPipe_ready;
  wire                readStage_controlPipe_payload_frameStart;
  wire                readStage_controlPipe_payload_rowEnd;
  wire                readStage_controlPipe_payload_pipeValid;
  wire                readStage_controlPipe_payload_firstRow;
  wire                readStage_controlPipe_payload_lastRow;
  wire                readStage_controlPipe_payload_finalResult;
  wire                readStage_controlPipe_payload_mainCompare;
  wire                readStage_controlPipe_payload_counterCompare;
  wire                readStage_controlPipe_payload_horizontalCompare;
  wire                readStage_controlPipe_payload_verticalCompare;
  wire       [7:0]    readStage_controlPipe_payload_mainDiff;
  wire       [7:0]    readStage_controlPipe_payload_counterDiff;
  wire       [7:0]    readStage_controlPipe_payload_horizontalDiff;
  wire       [7:0]    readStage_controlPipe_payload_verticalDiff;
  wire                readStage_controlPipe_payload_isHorizontalMin;
  wire       [7:0]    readStage_controlPipe_payload_minDiff;
  wire       [1:0]    readStage_controlPipe_payload_currentPosition;
  wire       [1:0]    readStage_controlPipe_payload_nextPosition;
  wire                readStage_controlPipe_payload_horizontalDirectionValid;
  wire                readStage_controlPipe_payload_verticalDirectionValid;
  wire                readStage_controlPipe_payload_mainDirectionValid;
  wire                readStage_controlPipe_payload_counterDirectionValid;
  wire                readStage_controlPipe_payload_inValidMinDiff;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_frameStart;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_rowEnd;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_pipeValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_firstRow;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_lastRow;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_finalResult;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainCompare;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterCompare;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_horizontalCompare;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_verticalCompare;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_horizontalDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_verticalDiff;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_isHorizontalMin;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_minDiff;
  reg        [1:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_currentPosition;
  reg        [1:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_nextPosition;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_horizontalDirectionValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_verticalDirectionValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainDirectionValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterDirectionValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_inValidMinDiff;
  wire                when_Stream_l368_27;
  wire                readStage_mainOnePixelStream_s2mPipe_valid;
  reg                 readStage_mainOnePixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_mainOnePixelStream_s2mPipe_payload;
  reg                 readStage_mainOnePixelStream_rValid;
  reg        [7:0]    readStage_mainOnePixelStream_rData;
  wire                compareStage_mainOnePixelStream_valid;
  wire                compareStage_mainOnePixelStream_ready;
  wire       [7:0]    compareStage_mainOnePixelStream_payload;
  reg                 readStage_mainOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_mainOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_28;
  wire                readStage_counterOnePixelStream_s2mPipe_valid;
  reg                 readStage_counterOnePixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_counterOnePixelStream_s2mPipe_payload;
  reg                 readStage_counterOnePixelStream_rValid;
  reg        [7:0]    readStage_counterOnePixelStream_rData;
  wire                compareStage_counterOnePixelStream_valid;
  wire                compareStage_counterOnePixelStream_ready;
  wire       [7:0]    compareStage_counterOnePixelStream_payload;
  reg                 readStage_counterOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_counterOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_29;
  wire                readStage_mainTwoPixelStream_s2mPipe_valid;
  reg                 readStage_mainTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_mainTwoPixelStream_s2mPipe_payload;
  reg                 readStage_mainTwoPixelStream_rValid;
  reg        [7:0]    readStage_mainTwoPixelStream_rData;
  wire                compareStage_mainTwoPixelStream_valid;
  wire                compareStage_mainTwoPixelStream_ready;
  wire       [7:0]    compareStage_mainTwoPixelStream_payload;
  reg                 readStage_mainTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_mainTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_30;
  wire                readStage_counterTwoPixelStream_s2mPipe_valid;
  reg                 readStage_counterTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_counterTwoPixelStream_s2mPipe_payload;
  reg                 readStage_counterTwoPixelStream_rValid;
  reg        [7:0]    readStage_counterTwoPixelStream_rData;
  wire                compareStage_counterTwoPixelStream_valid;
  wire                compareStage_counterTwoPixelStream_ready;
  wire       [7:0]    compareStage_counterTwoPixelStream_payload;
  reg                 readStage_counterTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_counterTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_31;
  wire                readStage_mainThreePixelStream_s2mPipe_valid;
  reg                 readStage_mainThreePixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_mainThreePixelStream_s2mPipe_payload;
  reg                 readStage_mainThreePixelStream_rValid;
  reg        [7:0]    readStage_mainThreePixelStream_rData;
  wire                compareStage_mainThreePixelStream_valid;
  wire                compareStage_mainThreePixelStream_ready;
  wire       [7:0]    compareStage_mainThreePixelStream_payload;
  reg                 readStage_mainThreePixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_mainThreePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_32;
  wire                readStage_counterThreePixelStream_s2mPipe_valid;
  reg                 readStage_counterThreePixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_counterThreePixelStream_s2mPipe_payload;
  reg                 readStage_counterThreePixelStream_rValid;
  reg        [7:0]    readStage_counterThreePixelStream_rData;
  wire                compareStage_counterThreePixelStream_valid;
  wire                compareStage_counterThreePixelStream_ready;
  wire       [7:0]    compareStage_counterThreePixelStream_payload;
  reg                 readStage_counterThreePixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_counterThreePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_33;
  wire                readStage_mainOneValidStream_s2mPipe_valid;
  reg                 readStage_mainOneValidStream_s2mPipe_ready;
  wire                readStage_mainOneValidStream_s2mPipe_payload;
  reg                 readStage_mainOneValidStream_rValid;
  reg                 readStage_mainOneValidStream_rData;
  wire                compareStage_mainOneValidStream_valid;
  wire                compareStage_mainOneValidStream_ready;
  wire                compareStage_mainOneValidStream_payload;
  reg                 readStage_mainOneValidStream_s2mPipe_rValid;
  reg                 readStage_mainOneValidStream_s2mPipe_rData;
  wire                when_Stream_l368_34;
  wire                readStage_counterOneValidStream_s2mPipe_valid;
  reg                 readStage_counterOneValidStream_s2mPipe_ready;
  wire                readStage_counterOneValidStream_s2mPipe_payload;
  reg                 readStage_counterOneValidStream_rValid;
  reg                 readStage_counterOneValidStream_rData;
  wire                compareStage_counterOneValidStream_valid;
  wire                compareStage_counterOneValidStream_ready;
  wire                compareStage_counterOneValidStream_payload;
  reg                 readStage_counterOneValidStream_s2mPipe_rValid;
  reg                 readStage_counterOneValidStream_s2mPipe_rData;
  wire                when_Stream_l368_35;
  wire                readStage_mainTwoValidStream_s2mPipe_valid;
  reg                 readStage_mainTwoValidStream_s2mPipe_ready;
  wire                readStage_mainTwoValidStream_s2mPipe_payload;
  reg                 readStage_mainTwoValidStream_rValid;
  reg                 readStage_mainTwoValidStream_rData;
  wire                compareStage_mainTwoValidStream_valid;
  wire                compareStage_mainTwoValidStream_ready;
  wire                compareStage_mainTwoValidStream_payload;
  reg                 readStage_mainTwoValidStream_s2mPipe_rValid;
  reg                 readStage_mainTwoValidStream_s2mPipe_rData;
  wire                when_Stream_l368_36;
  wire                readStage_counterTwoValidStream_s2mPipe_valid;
  reg                 readStage_counterTwoValidStream_s2mPipe_ready;
  wire                readStage_counterTwoValidStream_s2mPipe_payload;
  reg                 readStage_counterTwoValidStream_rValid;
  reg                 readStage_counterTwoValidStream_rData;
  wire                compareStage_counterTwoValidStream_valid;
  wire                compareStage_counterTwoValidStream_ready;
  wire                compareStage_counterTwoValidStream_payload;
  reg                 readStage_counterTwoValidStream_s2mPipe_rValid;
  reg                 readStage_counterTwoValidStream_s2mPipe_rData;
  wire                when_Stream_l368_37;
  wire                readStage_mainThreeValidStream_s2mPipe_valid;
  reg                 readStage_mainThreeValidStream_s2mPipe_ready;
  wire                readStage_mainThreeValidStream_s2mPipe_payload;
  reg                 readStage_mainThreeValidStream_rValid;
  reg                 readStage_mainThreeValidStream_rData;
  wire                compareStage_mainThreeValidStream_valid;
  wire                compareStage_mainThreeValidStream_ready;
  wire                compareStage_mainThreeValidStream_payload;
  reg                 readStage_mainThreeValidStream_s2mPipe_rValid;
  reg                 readStage_mainThreeValidStream_s2mPipe_rData;
  wire                when_Stream_l368_38;
  wire                readStage_counterThreeValidStream_s2mPipe_valid;
  reg                 readStage_counterThreeValidStream_s2mPipe_ready;
  wire                readStage_counterThreeValidStream_s2mPipe_payload;
  reg                 readStage_counterThreeValidStream_rValid;
  reg                 readStage_counterThreeValidStream_rData;
  wire                compareStage_counterThreeValidStream_valid;
  wire                compareStage_counterThreeValidStream_ready;
  wire                compareStage_counterThreeValidStream_payload;
  reg                 readStage_counterThreeValidStream_s2mPipe_rValid;
  reg                 readStage_counterThreeValidStream_s2mPipe_rData;
  wire                when_Stream_l368_39;
  reg                 CICC1851_readStage_controlPipe_translated_payload_mainCompare;
  reg                 CICC1851_readStage_controlPipe_translated_payload_counterCompare;
  reg                 CICC1851_readStage_controlPipe_translated_payload_horizontalCompare;
  reg                 CICC1851_readStage_controlPipe_translated_payload_verticalCompare;
  reg                 CICC1851_readStage_controlPipe_translated_payload_horizontalDirectionValid;
  reg                 CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid;
  reg                 CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid;
  reg                 CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid;
  wire                when_SuperResolutionPart3_l342;
  wire                when_SuperResolutionPart3_l344;
  wire                when_SuperResolutionPart3_l345;
  wire                when_SuperResolutionPart3_l348;
  wire                when_SuperResolutionPart3_l351;
  wire                when_SuperResolutionPart3_l347;
  wire                when_SuperResolutionPart3_l356;
  wire                when_SuperResolutionPart3_l357;
  wire                when_SuperResolutionPart3_l365;
  wire                when_SuperResolutionPart3_l373;
  wire                when_SuperResolutionPart3_l378;
  wire                when_SuperResolutionPart3_l383;
  wire                when_SuperResolutionPart3_l391;
  wire                when_SuperResolutionPart3_l396;
  wire                when_SuperResolutionPart3_l401;
  wire                when_SuperResolutionPart3_l409;
  wire                when_SuperResolutionPart3_l377;
  wire                when_SuperResolutionPart3_l415;
  wire                when_SuperResolutionPart3_l416;
  wire                when_SuperResolutionPart3_l419;
  wire                when_SuperResolutionPart3_l422;
  wire                when_SuperResolutionPart3_l424;
  wire                when_SuperResolutionPart3_l432;
  wire                when_SuperResolutionPart3_l441;
  wire                when_SuperResolutionPart3_l449;
  wire                when_SuperResolutionPart3_l458;
  wire                when_SuperResolutionPart3_l460;
  wire                when_SuperResolutionPart3_l463;
  wire                when_SuperResolutionPart3_l465;
  wire                when_SuperResolutionPart3_l470;
  wire                when_SuperResolutionPart3_l477;
  wire                when_SuperResolutionPart3_l485;
  wire                when_SuperResolutionPart3_l487;
  wire                when_SuperResolutionPart3_l490;
  wire                when_SuperResolutionPart3_l492;
  wire                when_SuperResolutionPart3_l497;
  wire                when_SuperResolutionPart3_l500;
  wire                when_SuperResolutionPart3_l502;
  wire                when_SuperResolutionPart3_l504;
  wire                when_SuperResolutionPart3_l511;
  wire                when_SuperResolutionPart3_l519;
  wire                when_SuperResolutionPart3_l521;
  wire                when_SuperResolutionPart3_l524;
  wire                when_SuperResolutionPart3_l526;
  wire                when_SuperResolutionPart3_l531;
  wire                when_SuperResolutionPart3_l539;
  wire                when_SuperResolutionPart3_l547;
  wire                when_SuperResolutionPart3_l549;
  wire                when_SuperResolutionPart3_l552;
  wire                when_SuperResolutionPart3_l554;
  wire                when_SuperResolutionPart3_l559;
  wire                when_SuperResolutionPart3_l562;
  wire                when_SuperResolutionPart3_l564;
  wire                when_SuperResolutionPart3_l566;
  wire                when_SuperResolutionPart3_l573;
  wire                when_SuperResolutionPart3_l581;
  wire                when_SuperResolutionPart3_l583;
  wire                when_SuperResolutionPart3_l586;
  wire                when_SuperResolutionPart3_l588;
  wire                when_SuperResolutionPart3_l593;
  wire                when_SuperResolutionPart3_l601;
  wire                when_SuperResolutionPart3_l609;
  wire                when_SuperResolutionPart3_l611;
  wire                when_SuperResolutionPart3_l614;
  wire                when_SuperResolutionPart3_l616;
  wire                when_SuperResolutionPart3_l496;
  wire                readStage_controlPipe_translated_valid;
  wire                readStage_controlPipe_translated_ready;
  wire                readStage_controlPipe_translated_payload_frameStart;
  wire                readStage_controlPipe_translated_payload_rowEnd;
  wire                readStage_controlPipe_translated_payload_pipeValid;
  wire                readStage_controlPipe_translated_payload_firstRow;
  wire                readStage_controlPipe_translated_payload_lastRow;
  wire                readStage_controlPipe_translated_payload_finalResult;
  wire                readStage_controlPipe_translated_payload_mainCompare;
  wire                readStage_controlPipe_translated_payload_counterCompare;
  wire                readStage_controlPipe_translated_payload_horizontalCompare;
  wire                readStage_controlPipe_translated_payload_verticalCompare;
  wire       [7:0]    readStage_controlPipe_translated_payload_mainDiff;
  wire       [7:0]    readStage_controlPipe_translated_payload_counterDiff;
  wire       [7:0]    readStage_controlPipe_translated_payload_horizontalDiff;
  wire       [7:0]    readStage_controlPipe_translated_payload_verticalDiff;
  wire                readStage_controlPipe_translated_payload_isHorizontalMin;
  wire       [7:0]    readStage_controlPipe_translated_payload_minDiff;
  wire       [1:0]    readStage_controlPipe_translated_payload_currentPosition;
  wire       [1:0]    readStage_controlPipe_translated_payload_nextPosition;
  wire                readStage_controlPipe_translated_payload_horizontalDirectionValid;
  wire                readStage_controlPipe_translated_payload_verticalDirectionValid;
  wire                readStage_controlPipe_translated_payload_mainDirectionValid;
  wire                readStage_controlPipe_translated_payload_counterDirectionValid;
  wire                readStage_controlPipe_translated_payload_inValidMinDiff;
  wire                readStage_controlPipe_translated_s2mPipe_valid;
  reg                 readStage_controlPipe_translated_s2mPipe_ready;
  wire                readStage_controlPipe_translated_s2mPipe_payload_frameStart;
  wire                readStage_controlPipe_translated_s2mPipe_payload_rowEnd;
  wire                readStage_controlPipe_translated_s2mPipe_payload_pipeValid;
  wire                readStage_controlPipe_translated_s2mPipe_payload_firstRow;
  wire                readStage_controlPipe_translated_s2mPipe_payload_lastRow;
  wire                readStage_controlPipe_translated_s2mPipe_payload_finalResult;
  wire                readStage_controlPipe_translated_s2mPipe_payload_mainCompare;
  wire                readStage_controlPipe_translated_s2mPipe_payload_counterCompare;
  wire                readStage_controlPipe_translated_s2mPipe_payload_horizontalCompare;
  wire                readStage_controlPipe_translated_s2mPipe_payload_verticalCompare;
  wire       [7:0]    readStage_controlPipe_translated_s2mPipe_payload_mainDiff;
  wire       [7:0]    readStage_controlPipe_translated_s2mPipe_payload_counterDiff;
  wire       [7:0]    readStage_controlPipe_translated_s2mPipe_payload_horizontalDiff;
  wire       [7:0]    readStage_controlPipe_translated_s2mPipe_payload_verticalDiff;
  wire                readStage_controlPipe_translated_s2mPipe_payload_isHorizontalMin;
  wire       [7:0]    readStage_controlPipe_translated_s2mPipe_payload_minDiff;
  wire       [1:0]    readStage_controlPipe_translated_s2mPipe_payload_currentPosition;
  wire       [1:0]    readStage_controlPipe_translated_s2mPipe_payload_nextPosition;
  wire                readStage_controlPipe_translated_s2mPipe_payload_horizontalDirectionValid;
  wire                readStage_controlPipe_translated_s2mPipe_payload_verticalDirectionValid;
  wire                readStage_controlPipe_translated_s2mPipe_payload_mainDirectionValid;
  wire                readStage_controlPipe_translated_s2mPipe_payload_counterDirectionValid;
  wire                readStage_controlPipe_translated_s2mPipe_payload_inValidMinDiff;
  reg                 readStage_controlPipe_translated_rValid;
  reg                 readStage_controlPipe_translated_rData_frameStart;
  reg                 readStage_controlPipe_translated_rData_rowEnd;
  reg                 readStage_controlPipe_translated_rData_pipeValid;
  reg                 readStage_controlPipe_translated_rData_firstRow;
  reg                 readStage_controlPipe_translated_rData_lastRow;
  reg                 readStage_controlPipe_translated_rData_finalResult;
  reg                 readStage_controlPipe_translated_rData_mainCompare;
  reg                 readStage_controlPipe_translated_rData_counterCompare;
  reg                 readStage_controlPipe_translated_rData_horizontalCompare;
  reg                 readStage_controlPipe_translated_rData_verticalCompare;
  reg        [7:0]    readStage_controlPipe_translated_rData_mainDiff;
  reg        [7:0]    readStage_controlPipe_translated_rData_counterDiff;
  reg        [7:0]    readStage_controlPipe_translated_rData_horizontalDiff;
  reg        [7:0]    readStage_controlPipe_translated_rData_verticalDiff;
  reg                 readStage_controlPipe_translated_rData_isHorizontalMin;
  reg        [7:0]    readStage_controlPipe_translated_rData_minDiff;
  reg        [1:0]    readStage_controlPipe_translated_rData_currentPosition;
  reg        [1:0]    readStage_controlPipe_translated_rData_nextPosition;
  reg                 readStage_controlPipe_translated_rData_horizontalDirectionValid;
  reg                 readStage_controlPipe_translated_rData_verticalDirectionValid;
  reg                 readStage_controlPipe_translated_rData_mainDirectionValid;
  reg                 readStage_controlPipe_translated_rData_counterDirectionValid;
  reg                 readStage_controlPipe_translated_rData_inValidMinDiff;
  wire                compareStage_controlPipe_valid;
  wire                compareStage_controlPipe_ready;
  wire                compareStage_controlPipe_payload_frameStart;
  wire                compareStage_controlPipe_payload_rowEnd;
  wire                compareStage_controlPipe_payload_pipeValid;
  wire                compareStage_controlPipe_payload_firstRow;
  wire                compareStage_controlPipe_payload_lastRow;
  wire                compareStage_controlPipe_payload_finalResult;
  wire                compareStage_controlPipe_payload_mainCompare;
  wire                compareStage_controlPipe_payload_counterCompare;
  wire                compareStage_controlPipe_payload_horizontalCompare;
  wire                compareStage_controlPipe_payload_verticalCompare;
  wire       [7:0]    compareStage_controlPipe_payload_mainDiff;
  wire       [7:0]    compareStage_controlPipe_payload_counterDiff;
  wire       [7:0]    compareStage_controlPipe_payload_horizontalDiff;
  wire       [7:0]    compareStage_controlPipe_payload_verticalDiff;
  wire                compareStage_controlPipe_payload_isHorizontalMin;
  wire       [7:0]    compareStage_controlPipe_payload_minDiff;
  wire       [1:0]    compareStage_controlPipe_payload_currentPosition;
  wire       [1:0]    compareStage_controlPipe_payload_nextPosition;
  wire                compareStage_controlPipe_payload_horizontalDirectionValid;
  wire                compareStage_controlPipe_payload_verticalDirectionValid;
  wire                compareStage_controlPipe_payload_mainDirectionValid;
  wire                compareStage_controlPipe_payload_counterDirectionValid;
  wire                compareStage_controlPipe_payload_inValidMinDiff;
  reg                 readStage_controlPipe_translated_s2mPipe_rValid;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_frameStart;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_rowEnd;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_pipeValid;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_firstRow;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_lastRow;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_finalResult;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_mainCompare;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_counterCompare;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_horizontalCompare;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_verticalCompare;
  reg        [7:0]    readStage_controlPipe_translated_s2mPipe_rData_mainDiff;
  reg        [7:0]    readStage_controlPipe_translated_s2mPipe_rData_counterDiff;
  reg        [7:0]    readStage_controlPipe_translated_s2mPipe_rData_horizontalDiff;
  reg        [7:0]    readStage_controlPipe_translated_s2mPipe_rData_verticalDiff;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_isHorizontalMin;
  reg        [7:0]    readStage_controlPipe_translated_s2mPipe_rData_minDiff;
  reg        [1:0]    readStage_controlPipe_translated_s2mPipe_rData_currentPosition;
  reg        [1:0]    readStage_controlPipe_translated_s2mPipe_rData_nextPosition;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_horizontalDirectionValid;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_verticalDirectionValid;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_mainDirectionValid;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_counterDirectionValid;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_inValidMinDiff;
  wire                when_Stream_l368_40;
  wire                compareStage_mainOnePixelStream_s2mPipe_valid;
  reg                 compareStage_mainOnePixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_mainOnePixelStream_s2mPipe_payload;
  reg                 compareStage_mainOnePixelStream_rValid;
  reg        [7:0]    compareStage_mainOnePixelStream_rData;
  wire                diffStage_mainOnePixelStream_valid;
  wire                diffStage_mainOnePixelStream_ready;
  wire       [7:0]    diffStage_mainOnePixelStream_payload;
  reg                 compareStage_mainOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_mainOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_41;
  wire                compareStage_counterOnePixelStream_s2mPipe_valid;
  reg                 compareStage_counterOnePixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_counterOnePixelStream_s2mPipe_payload;
  reg                 compareStage_counterOnePixelStream_rValid;
  reg        [7:0]    compareStage_counterOnePixelStream_rData;
  wire                diffStage_counterOnePixelStream_valid;
  wire                diffStage_counterOnePixelStream_ready;
  wire       [7:0]    diffStage_counterOnePixelStream_payload;
  reg                 compareStage_counterOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_counterOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_42;
  wire                compareStage_mainTwoPixelStream_s2mPipe_valid;
  reg                 compareStage_mainTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_mainTwoPixelStream_s2mPipe_payload;
  reg                 compareStage_mainTwoPixelStream_rValid;
  reg        [7:0]    compareStage_mainTwoPixelStream_rData;
  wire                diffStage_mainTwoPixelStream_valid;
  wire                diffStage_mainTwoPixelStream_ready;
  wire       [7:0]    diffStage_mainTwoPixelStream_payload;
  reg                 compareStage_mainTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_mainTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_43;
  wire                compareStage_counterTwoPixelStream_s2mPipe_valid;
  reg                 compareStage_counterTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_counterTwoPixelStream_s2mPipe_payload;
  reg                 compareStage_counterTwoPixelStream_rValid;
  reg        [7:0]    compareStage_counterTwoPixelStream_rData;
  wire                diffStage_counterTwoPixelStream_valid;
  wire                diffStage_counterTwoPixelStream_ready;
  wire       [7:0]    diffStage_counterTwoPixelStream_payload;
  reg                 compareStage_counterTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_counterTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_44;
  wire                compareStage_mainThreePixelStream_s2mPipe_valid;
  reg                 compareStage_mainThreePixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_mainThreePixelStream_s2mPipe_payload;
  reg                 compareStage_mainThreePixelStream_rValid;
  reg        [7:0]    compareStage_mainThreePixelStream_rData;
  wire                diffStage_mainThreePixelStream_valid;
  wire                diffStage_mainThreePixelStream_ready;
  wire       [7:0]    diffStage_mainThreePixelStream_payload;
  reg                 compareStage_mainThreePixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_mainThreePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_45;
  wire                compareStage_counterThreePixelStream_s2mPipe_valid;
  reg                 compareStage_counterThreePixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_counterThreePixelStream_s2mPipe_payload;
  reg                 compareStage_counterThreePixelStream_rValid;
  reg        [7:0]    compareStage_counterThreePixelStream_rData;
  wire                diffStage_counterThreePixelStream_valid;
  wire                diffStage_counterThreePixelStream_ready;
  wire       [7:0]    diffStage_counterThreePixelStream_payload;
  reg                 compareStage_counterThreePixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_counterThreePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_46;
  wire                compareStage_mainOneValidStream_s2mPipe_valid;
  reg                 compareStage_mainOneValidStream_s2mPipe_ready;
  wire                compareStage_mainOneValidStream_s2mPipe_payload;
  reg                 compareStage_mainOneValidStream_rValid;
  reg                 compareStage_mainOneValidStream_rData;
  wire                diffStage_mainOneValidStream_valid;
  wire                diffStage_mainOneValidStream_ready;
  wire                diffStage_mainOneValidStream_payload;
  reg                 compareStage_mainOneValidStream_s2mPipe_rValid;
  reg                 compareStage_mainOneValidStream_s2mPipe_rData;
  wire                when_Stream_l368_47;
  wire                compareStage_counterOneValidStream_s2mPipe_valid;
  reg                 compareStage_counterOneValidStream_s2mPipe_ready;
  wire                compareStage_counterOneValidStream_s2mPipe_payload;
  reg                 compareStage_counterOneValidStream_rValid;
  reg                 compareStage_counterOneValidStream_rData;
  wire                diffStage_counterOneValidStream_valid;
  wire                diffStage_counterOneValidStream_ready;
  wire                diffStage_counterOneValidStream_payload;
  reg                 compareStage_counterOneValidStream_s2mPipe_rValid;
  reg                 compareStage_counterOneValidStream_s2mPipe_rData;
  wire                when_Stream_l368_48;
  wire                compareStage_mainTwoValidStream_s2mPipe_valid;
  reg                 compareStage_mainTwoValidStream_s2mPipe_ready;
  wire                compareStage_mainTwoValidStream_s2mPipe_payload;
  reg                 compareStage_mainTwoValidStream_rValid;
  reg                 compareStage_mainTwoValidStream_rData;
  wire                diffStage_mainTwoValidStream_valid;
  wire                diffStage_mainTwoValidStream_ready;
  wire                diffStage_mainTwoValidStream_payload;
  reg                 compareStage_mainTwoValidStream_s2mPipe_rValid;
  reg                 compareStage_mainTwoValidStream_s2mPipe_rData;
  wire                when_Stream_l368_49;
  wire                compareStage_counterTwoValidStream_s2mPipe_valid;
  reg                 compareStage_counterTwoValidStream_s2mPipe_ready;
  wire                compareStage_counterTwoValidStream_s2mPipe_payload;
  reg                 compareStage_counterTwoValidStream_rValid;
  reg                 compareStage_counterTwoValidStream_rData;
  wire                diffStage_counterTwoValidStream_valid;
  wire                diffStage_counterTwoValidStream_ready;
  wire                diffStage_counterTwoValidStream_payload;
  reg                 compareStage_counterTwoValidStream_s2mPipe_rValid;
  reg                 compareStage_counterTwoValidStream_s2mPipe_rData;
  wire                when_Stream_l368_50;
  wire                compareStage_mainThreeValidStream_s2mPipe_valid;
  reg                 compareStage_mainThreeValidStream_s2mPipe_ready;
  wire                compareStage_mainThreeValidStream_s2mPipe_payload;
  reg                 compareStage_mainThreeValidStream_rValid;
  reg                 compareStage_mainThreeValidStream_rData;
  wire                diffStage_mainThreeValidStream_valid;
  wire                diffStage_mainThreeValidStream_ready;
  wire                diffStage_mainThreeValidStream_payload;
  reg                 compareStage_mainThreeValidStream_s2mPipe_rValid;
  reg                 compareStage_mainThreeValidStream_s2mPipe_rData;
  wire                when_Stream_l368_51;
  wire                compareStage_counterThreeValidStream_s2mPipe_valid;
  reg                 compareStage_counterThreeValidStream_s2mPipe_ready;
  wire                compareStage_counterThreeValidStream_s2mPipe_payload;
  reg                 compareStage_counterThreeValidStream_rValid;
  reg                 compareStage_counterThreeValidStream_rData;
  wire                diffStage_counterThreeValidStream_valid;
  wire                diffStage_counterThreeValidStream_ready;
  wire                diffStage_counterThreeValidStream_payload;
  reg                 compareStage_counterThreeValidStream_s2mPipe_rValid;
  reg                 compareStage_counterThreeValidStream_s2mPipe_rData;
  wire                when_Stream_l368_52;
  reg        [7:0]    CICC1851_compareStage_controlPipe_translated_payload_mainDiff;
  reg        [7:0]    CICC1851_compareStage_controlPipe_translated_payload_counterDiff;
  reg        [7:0]    CICC1851_compareStage_controlPipe_translated_payload_horizontalDiff;
  reg        [7:0]    CICC1851_compareStage_controlPipe_translated_payload_verticalDiff;
  reg                 CICC1851_compareStage_controlPipe_translated_payload_inValidMinDiff;
  wire                when_SuperResolutionPart3_l647;
  wire                when_SuperResolutionPart3_l649;
  wire                when_SuperResolutionPart3_l652;
  wire                when_SuperResolutionPart3_l661;
  wire                when_SuperResolutionPart3_l664;
  wire                when_SuperResolutionPart3_l697;
  wire                when_SuperResolutionPart3_l725;
  wire                when_SuperResolutionPart3_l694;
  wire                when_SuperResolutionPart3_l753;
  wire                compareStage_controlPipe_translated_valid;
  wire                compareStage_controlPipe_translated_ready;
  wire                compareStage_controlPipe_translated_payload_frameStart;
  wire                compareStage_controlPipe_translated_payload_rowEnd;
  wire                compareStage_controlPipe_translated_payload_pipeValid;
  wire                compareStage_controlPipe_translated_payload_firstRow;
  wire                compareStage_controlPipe_translated_payload_lastRow;
  wire                compareStage_controlPipe_translated_payload_finalResult;
  wire                compareStage_controlPipe_translated_payload_mainCompare;
  wire                compareStage_controlPipe_translated_payload_counterCompare;
  wire                compareStage_controlPipe_translated_payload_horizontalCompare;
  wire                compareStage_controlPipe_translated_payload_verticalCompare;
  wire       [7:0]    compareStage_controlPipe_translated_payload_mainDiff;
  wire       [7:0]    compareStage_controlPipe_translated_payload_counterDiff;
  wire       [7:0]    compareStage_controlPipe_translated_payload_horizontalDiff;
  wire       [7:0]    compareStage_controlPipe_translated_payload_verticalDiff;
  wire                compareStage_controlPipe_translated_payload_isHorizontalMin;
  wire       [7:0]    compareStage_controlPipe_translated_payload_minDiff;
  wire       [1:0]    compareStage_controlPipe_translated_payload_currentPosition;
  wire       [1:0]    compareStage_controlPipe_translated_payload_nextPosition;
  wire                compareStage_controlPipe_translated_payload_horizontalDirectionValid;
  wire                compareStage_controlPipe_translated_payload_verticalDirectionValid;
  wire                compareStage_controlPipe_translated_payload_mainDirectionValid;
  wire                compareStage_controlPipe_translated_payload_counterDirectionValid;
  wire                compareStage_controlPipe_translated_payload_inValidMinDiff;
  wire                compareStage_controlPipe_translated_s2mPipe_valid;
  reg                 compareStage_controlPipe_translated_s2mPipe_ready;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_frameStart;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_rowEnd;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_pipeValid;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_firstRow;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_lastRow;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_finalResult;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_mainCompare;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_counterCompare;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_horizontalCompare;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_verticalCompare;
  wire       [7:0]    compareStage_controlPipe_translated_s2mPipe_payload_mainDiff;
  wire       [7:0]    compareStage_controlPipe_translated_s2mPipe_payload_counterDiff;
  wire       [7:0]    compareStage_controlPipe_translated_s2mPipe_payload_horizontalDiff;
  wire       [7:0]    compareStage_controlPipe_translated_s2mPipe_payload_verticalDiff;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_isHorizontalMin;
  wire       [7:0]    compareStage_controlPipe_translated_s2mPipe_payload_minDiff;
  wire       [1:0]    compareStage_controlPipe_translated_s2mPipe_payload_currentPosition;
  wire       [1:0]    compareStage_controlPipe_translated_s2mPipe_payload_nextPosition;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_horizontalDirectionValid;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_verticalDirectionValid;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_mainDirectionValid;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_counterDirectionValid;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_inValidMinDiff;
  reg                 compareStage_controlPipe_translated_rValid;
  reg                 compareStage_controlPipe_translated_rData_frameStart;
  reg                 compareStage_controlPipe_translated_rData_rowEnd;
  reg                 compareStage_controlPipe_translated_rData_pipeValid;
  reg                 compareStage_controlPipe_translated_rData_firstRow;
  reg                 compareStage_controlPipe_translated_rData_lastRow;
  reg                 compareStage_controlPipe_translated_rData_finalResult;
  reg                 compareStage_controlPipe_translated_rData_mainCompare;
  reg                 compareStage_controlPipe_translated_rData_counterCompare;
  reg                 compareStage_controlPipe_translated_rData_horizontalCompare;
  reg                 compareStage_controlPipe_translated_rData_verticalCompare;
  reg        [7:0]    compareStage_controlPipe_translated_rData_mainDiff;
  reg        [7:0]    compareStage_controlPipe_translated_rData_counterDiff;
  reg        [7:0]    compareStage_controlPipe_translated_rData_horizontalDiff;
  reg        [7:0]    compareStage_controlPipe_translated_rData_verticalDiff;
  reg                 compareStage_controlPipe_translated_rData_isHorizontalMin;
  reg        [7:0]    compareStage_controlPipe_translated_rData_minDiff;
  reg        [1:0]    compareStage_controlPipe_translated_rData_currentPosition;
  reg        [1:0]    compareStage_controlPipe_translated_rData_nextPosition;
  reg                 compareStage_controlPipe_translated_rData_horizontalDirectionValid;
  reg                 compareStage_controlPipe_translated_rData_verticalDirectionValid;
  reg                 compareStage_controlPipe_translated_rData_mainDirectionValid;
  reg                 compareStage_controlPipe_translated_rData_counterDirectionValid;
  reg                 compareStage_controlPipe_translated_rData_inValidMinDiff;
  wire                diffStage_controlPipe_valid;
  wire                diffStage_controlPipe_ready;
  wire                diffStage_controlPipe_payload_frameStart;
  wire                diffStage_controlPipe_payload_rowEnd;
  wire                diffStage_controlPipe_payload_pipeValid;
  wire                diffStage_controlPipe_payload_firstRow;
  wire                diffStage_controlPipe_payload_lastRow;
  wire                diffStage_controlPipe_payload_finalResult;
  wire                diffStage_controlPipe_payload_mainCompare;
  wire                diffStage_controlPipe_payload_counterCompare;
  wire                diffStage_controlPipe_payload_horizontalCompare;
  wire                diffStage_controlPipe_payload_verticalCompare;
  wire       [7:0]    diffStage_controlPipe_payload_mainDiff;
  wire       [7:0]    diffStage_controlPipe_payload_counterDiff;
  wire       [7:0]    diffStage_controlPipe_payload_horizontalDiff;
  wire       [7:0]    diffStage_controlPipe_payload_verticalDiff;
  wire                diffStage_controlPipe_payload_isHorizontalMin;
  wire       [7:0]    diffStage_controlPipe_payload_minDiff;
  wire       [1:0]    diffStage_controlPipe_payload_currentPosition;
  wire       [1:0]    diffStage_controlPipe_payload_nextPosition;
  wire                diffStage_controlPipe_payload_horizontalDirectionValid;
  wire                diffStage_controlPipe_payload_verticalDirectionValid;
  wire                diffStage_controlPipe_payload_mainDirectionValid;
  wire                diffStage_controlPipe_payload_counterDirectionValid;
  wire                diffStage_controlPipe_payload_inValidMinDiff;
  reg                 compareStage_controlPipe_translated_s2mPipe_rValid;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_frameStart;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_rowEnd;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_pipeValid;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_firstRow;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_lastRow;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_finalResult;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_mainCompare;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_counterCompare;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_horizontalCompare;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_verticalCompare;
  reg        [7:0]    compareStage_controlPipe_translated_s2mPipe_rData_mainDiff;
  reg        [7:0]    compareStage_controlPipe_translated_s2mPipe_rData_counterDiff;
  reg        [7:0]    compareStage_controlPipe_translated_s2mPipe_rData_horizontalDiff;
  reg        [7:0]    compareStage_controlPipe_translated_s2mPipe_rData_verticalDiff;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_isHorizontalMin;
  reg        [7:0]    compareStage_controlPipe_translated_s2mPipe_rData_minDiff;
  reg        [1:0]    compareStage_controlPipe_translated_s2mPipe_rData_currentPosition;
  reg        [1:0]    compareStage_controlPipe_translated_s2mPipe_rData_nextPosition;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_horizontalDirectionValid;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_verticalDirectionValid;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_mainDirectionValid;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_counterDirectionValid;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_inValidMinDiff;
  wire                when_Stream_l368_53;
  wire                diffStage_mainOnePixelStream_s2mPipe_valid;
  reg                 diffStage_mainOnePixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_mainOnePixelStream_s2mPipe_payload;
  reg                 diffStage_mainOnePixelStream_rValid;
  reg        [7:0]    diffStage_mainOnePixelStream_rData;
  wire                resultStage_mainOnePixelStream_valid;
  wire                resultStage_mainOnePixelStream_ready;
  wire       [7:0]    resultStage_mainOnePixelStream_payload;
  reg                 diffStage_mainOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_mainOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_54;
  wire                diffStage_counterOnePixelStream_s2mPipe_valid;
  reg                 diffStage_counterOnePixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_counterOnePixelStream_s2mPipe_payload;
  reg                 diffStage_counterOnePixelStream_rValid;
  reg        [7:0]    diffStage_counterOnePixelStream_rData;
  wire                resultStage_counterOnePixelStream_valid;
  wire                resultStage_counterOnePixelStream_ready;
  wire       [7:0]    resultStage_counterOnePixelStream_payload;
  reg                 diffStage_counterOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_counterOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_55;
  wire                diffStage_mainTwoPixelStream_s2mPipe_valid;
  reg                 diffStage_mainTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_mainTwoPixelStream_s2mPipe_payload;
  reg                 diffStage_mainTwoPixelStream_rValid;
  reg        [7:0]    diffStage_mainTwoPixelStream_rData;
  wire                resultStage_mainTwoPixelStream_valid;
  wire                resultStage_mainTwoPixelStream_ready;
  wire       [7:0]    resultStage_mainTwoPixelStream_payload;
  reg                 diffStage_mainTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_mainTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_56;
  wire                diffStage_counterTwoPixelStream_s2mPipe_valid;
  reg                 diffStage_counterTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_counterTwoPixelStream_s2mPipe_payload;
  reg                 diffStage_counterTwoPixelStream_rValid;
  reg        [7:0]    diffStage_counterTwoPixelStream_rData;
  wire                resultStage_counterTwoPixelStream_valid;
  wire                resultStage_counterTwoPixelStream_ready;
  wire       [7:0]    resultStage_counterTwoPixelStream_payload;
  reg                 diffStage_counterTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_counterTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_57;
  wire                diffStage_mainThreePixelStream_s2mPipe_valid;
  reg                 diffStage_mainThreePixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_mainThreePixelStream_s2mPipe_payload;
  reg                 diffStage_mainThreePixelStream_rValid;
  reg        [7:0]    diffStage_mainThreePixelStream_rData;
  wire                resultStage_mainThreePixelStream_valid;
  wire                resultStage_mainThreePixelStream_ready;
  wire       [7:0]    resultStage_mainThreePixelStream_payload;
  reg                 diffStage_mainThreePixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_mainThreePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_58;
  wire                diffStage_counterThreePixelStream_s2mPipe_valid;
  reg                 diffStage_counterThreePixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_counterThreePixelStream_s2mPipe_payload;
  reg                 diffStage_counterThreePixelStream_rValid;
  reg        [7:0]    diffStage_counterThreePixelStream_rData;
  wire                resultStage_counterThreePixelStream_valid;
  wire                resultStage_counterThreePixelStream_ready;
  wire       [7:0]    resultStage_counterThreePixelStream_payload;
  reg                 diffStage_counterThreePixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_counterThreePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_59;
  wire                diffStage_mainOneValidStream_s2mPipe_valid;
  reg                 diffStage_mainOneValidStream_s2mPipe_ready;
  wire                diffStage_mainOneValidStream_s2mPipe_payload;
  reg                 diffStage_mainOneValidStream_rValid;
  reg                 diffStage_mainOneValidStream_rData;
  wire                resultStage_mainOneValidStream_valid;
  wire                resultStage_mainOneValidStream_ready;
  wire                resultStage_mainOneValidStream_payload;
  reg                 diffStage_mainOneValidStream_s2mPipe_rValid;
  reg                 diffStage_mainOneValidStream_s2mPipe_rData;
  wire                when_Stream_l368_60;
  wire                diffStage_counterOneValidStream_s2mPipe_valid;
  reg                 diffStage_counterOneValidStream_s2mPipe_ready;
  wire                diffStage_counterOneValidStream_s2mPipe_payload;
  reg                 diffStage_counterOneValidStream_rValid;
  reg                 diffStage_counterOneValidStream_rData;
  wire                resultStage_counterOneValidStream_valid;
  wire                resultStage_counterOneValidStream_ready;
  wire                resultStage_counterOneValidStream_payload;
  reg                 diffStage_counterOneValidStream_s2mPipe_rValid;
  reg                 diffStage_counterOneValidStream_s2mPipe_rData;
  wire                when_Stream_l368_61;
  wire                diffStage_mainTwoValidStream_s2mPipe_valid;
  reg                 diffStage_mainTwoValidStream_s2mPipe_ready;
  wire                diffStage_mainTwoValidStream_s2mPipe_payload;
  reg                 diffStage_mainTwoValidStream_rValid;
  reg                 diffStage_mainTwoValidStream_rData;
  wire                resultStage_mainTwoValidStream_valid;
  wire                resultStage_mainTwoValidStream_ready;
  wire                resultStage_mainTwoValidStream_payload;
  reg                 diffStage_mainTwoValidStream_s2mPipe_rValid;
  reg                 diffStage_mainTwoValidStream_s2mPipe_rData;
  wire                when_Stream_l368_62;
  wire                diffStage_counterTwoValidStream_s2mPipe_valid;
  reg                 diffStage_counterTwoValidStream_s2mPipe_ready;
  wire                diffStage_counterTwoValidStream_s2mPipe_payload;
  reg                 diffStage_counterTwoValidStream_rValid;
  reg                 diffStage_counterTwoValidStream_rData;
  wire                resultStage_counterTwoValidStream_valid;
  wire                resultStage_counterTwoValidStream_ready;
  wire                resultStage_counterTwoValidStream_payload;
  reg                 diffStage_counterTwoValidStream_s2mPipe_rValid;
  reg                 diffStage_counterTwoValidStream_s2mPipe_rData;
  wire                when_Stream_l368_63;
  wire                diffStage_mainThreeValidStream_s2mPipe_valid;
  reg                 diffStage_mainThreeValidStream_s2mPipe_ready;
  wire                diffStage_mainThreeValidStream_s2mPipe_payload;
  reg                 diffStage_mainThreeValidStream_rValid;
  reg                 diffStage_mainThreeValidStream_rData;
  wire                resultStage_mainThreeValidStream_valid;
  wire                resultStage_mainThreeValidStream_ready;
  wire                resultStage_mainThreeValidStream_payload;
  reg                 diffStage_mainThreeValidStream_s2mPipe_rValid;
  reg                 diffStage_mainThreeValidStream_s2mPipe_rData;
  wire                when_Stream_l368_64;
  wire                diffStage_counterThreeValidStream_s2mPipe_valid;
  reg                 diffStage_counterThreeValidStream_s2mPipe_ready;
  wire                diffStage_counterThreeValidStream_s2mPipe_payload;
  reg                 diffStage_counterThreeValidStream_rValid;
  reg                 diffStage_counterThreeValidStream_rData;
  wire                resultStage_counterThreeValidStream_valid;
  wire                resultStage_counterThreeValidStream_ready;
  wire                resultStage_counterThreeValidStream_payload;
  reg                 diffStage_counterThreeValidStream_s2mPipe_rValid;
  reg                 diffStage_counterThreeValidStream_s2mPipe_rData;
  wire                when_Stream_l368_65;
  reg                 CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin;
  reg        [7:0]    CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff;
  wire                when_SuperResolutionPart3_l783;
  wire                when_SuperResolutionPart3_l784;
  wire                when_SuperResolutionPart3_l785;
  wire                when_SuperResolutionPart3_l788;
  wire                when_SuperResolutionPart3_l796;
  wire                when_SuperResolutionPart3_l804;
  wire                when_SuperResolutionPart3_l812;
  wire                when_SuperResolutionPart3_l795;
  wire                when_SuperResolutionPart3_l803;
  wire                when_SuperResolutionPart3_l811;
  wire                when_SuperResolutionPart3_l819;
  wire                when_SuperResolutionPart3_l822;
  wire                when_SuperResolutionPart3_l825;
  wire                resultStage_controlPipeBeforePipe_valid;
  wire                resultStage_controlPipeBeforePipe_ready;
  wire                resultStage_controlPipeBeforePipe_payload_frameStart;
  wire                resultStage_controlPipeBeforePipe_payload_rowEnd;
  wire                resultStage_controlPipeBeforePipe_payload_pipeValid;
  wire                resultStage_controlPipeBeforePipe_payload_firstRow;
  wire                resultStage_controlPipeBeforePipe_payload_lastRow;
  wire                resultStage_controlPipeBeforePipe_payload_finalResult;
  wire                resultStage_controlPipeBeforePipe_payload_mainCompare;
  wire                resultStage_controlPipeBeforePipe_payload_counterCompare;
  wire                resultStage_controlPipeBeforePipe_payload_horizontalCompare;
  wire                resultStage_controlPipeBeforePipe_payload_verticalCompare;
  wire       [7:0]    resultStage_controlPipeBeforePipe_payload_mainDiff;
  wire       [7:0]    resultStage_controlPipeBeforePipe_payload_counterDiff;
  wire       [7:0]    resultStage_controlPipeBeforePipe_payload_horizontalDiff;
  wire       [7:0]    resultStage_controlPipeBeforePipe_payload_verticalDiff;
  wire                resultStage_controlPipeBeforePipe_payload_isHorizontalMin;
  wire       [7:0]    resultStage_controlPipeBeforePipe_payload_minDiff;
  wire       [1:0]    resultStage_controlPipeBeforePipe_payload_currentPosition;
  wire       [1:0]    resultStage_controlPipeBeforePipe_payload_nextPosition;
  wire                resultStage_controlPipeBeforePipe_payload_horizontalDirectionValid;
  wire                resultStage_controlPipeBeforePipe_payload_verticalDirectionValid;
  wire                resultStage_controlPipeBeforePipe_payload_mainDirectionValid;
  wire                resultStage_controlPipeBeforePipe_payload_counterDirectionValid;
  wire                resultStage_controlPipeBeforePipe_payload_inValidMinDiff;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_valid;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_ready;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_frameStart;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_rowEnd;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_pipeValid;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_firstRow;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_lastRow;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_finalResult;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_mainCompare;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_counterCompare;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_horizontalCompare;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_verticalCompare;
  wire       [7:0]    resultStage_controlPipeBeforePipe_s2mPipe_payload_mainDiff;
  wire       [7:0]    resultStage_controlPipeBeforePipe_s2mPipe_payload_counterDiff;
  wire       [7:0]    resultStage_controlPipeBeforePipe_s2mPipe_payload_horizontalDiff;
  wire       [7:0]    resultStage_controlPipeBeforePipe_s2mPipe_payload_verticalDiff;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_isHorizontalMin;
  wire       [7:0]    resultStage_controlPipeBeforePipe_s2mPipe_payload_minDiff;
  wire       [1:0]    resultStage_controlPipeBeforePipe_s2mPipe_payload_currentPosition;
  wire       [1:0]    resultStage_controlPipeBeforePipe_s2mPipe_payload_nextPosition;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_horizontalDirectionValid;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_verticalDirectionValid;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_mainDirectionValid;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_counterDirectionValid;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_inValidMinDiff;
  reg                 resultStage_controlPipeBeforePipe_rValid;
  reg                 resultStage_controlPipeBeforePipe_rData_frameStart;
  reg                 resultStage_controlPipeBeforePipe_rData_rowEnd;
  reg                 resultStage_controlPipeBeforePipe_rData_pipeValid;
  reg                 resultStage_controlPipeBeforePipe_rData_firstRow;
  reg                 resultStage_controlPipeBeforePipe_rData_lastRow;
  reg                 resultStage_controlPipeBeforePipe_rData_finalResult;
  reg                 resultStage_controlPipeBeforePipe_rData_mainCompare;
  reg                 resultStage_controlPipeBeforePipe_rData_counterCompare;
  reg                 resultStage_controlPipeBeforePipe_rData_horizontalCompare;
  reg                 resultStage_controlPipeBeforePipe_rData_verticalCompare;
  reg        [7:0]    resultStage_controlPipeBeforePipe_rData_mainDiff;
  reg        [7:0]    resultStage_controlPipeBeforePipe_rData_counterDiff;
  reg        [7:0]    resultStage_controlPipeBeforePipe_rData_horizontalDiff;
  reg        [7:0]    resultStage_controlPipeBeforePipe_rData_verticalDiff;
  reg                 resultStage_controlPipeBeforePipe_rData_isHorizontalMin;
  reg        [7:0]    resultStage_controlPipeBeforePipe_rData_minDiff;
  reg        [1:0]    resultStage_controlPipeBeforePipe_rData_currentPosition;
  reg        [1:0]    resultStage_controlPipeBeforePipe_rData_nextPosition;
  reg                 resultStage_controlPipeBeforePipe_rData_horizontalDirectionValid;
  reg                 resultStage_controlPipeBeforePipe_rData_verticalDirectionValid;
  reg                 resultStage_controlPipeBeforePipe_rData_mainDirectionValid;
  reg                 resultStage_controlPipeBeforePipe_rData_counterDirectionValid;
  reg                 resultStage_controlPipeBeforePipe_rData_inValidMinDiff;
  wire                resultStage_controlPipe_valid;
  wire                resultStage_controlPipe_ready;
  wire                resultStage_controlPipe_payload_frameStart;
  wire                resultStage_controlPipe_payload_rowEnd;
  wire                resultStage_controlPipe_payload_pipeValid;
  wire                resultStage_controlPipe_payload_firstRow;
  wire                resultStage_controlPipe_payload_lastRow;
  wire                resultStage_controlPipe_payload_finalResult;
  wire                resultStage_controlPipe_payload_mainCompare;
  wire                resultStage_controlPipe_payload_counterCompare;
  wire                resultStage_controlPipe_payload_horizontalCompare;
  wire                resultStage_controlPipe_payload_verticalCompare;
  wire       [7:0]    resultStage_controlPipe_payload_mainDiff;
  wire       [7:0]    resultStage_controlPipe_payload_counterDiff;
  wire       [7:0]    resultStage_controlPipe_payload_horizontalDiff;
  wire       [7:0]    resultStage_controlPipe_payload_verticalDiff;
  wire                resultStage_controlPipe_payload_isHorizontalMin;
  wire       [7:0]    resultStage_controlPipe_payload_minDiff;
  wire       [1:0]    resultStage_controlPipe_payload_currentPosition;
  wire       [1:0]    resultStage_controlPipe_payload_nextPosition;
  wire                resultStage_controlPipe_payload_horizontalDirectionValid;
  wire                resultStage_controlPipe_payload_verticalDirectionValid;
  wire                resultStage_controlPipe_payload_mainDirectionValid;
  wire                resultStage_controlPipe_payload_counterDirectionValid;
  wire                resultStage_controlPipe_payload_inValidMinDiff;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rValid;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_frameStart;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_rowEnd;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_pipeValid;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_firstRow;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_lastRow;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_finalResult;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_mainCompare;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_counterCompare;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_horizontalCompare;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_verticalCompare;
  reg        [7:0]    resultStage_controlPipeBeforePipe_s2mPipe_rData_mainDiff;
  reg        [7:0]    resultStage_controlPipeBeforePipe_s2mPipe_rData_counterDiff;
  reg        [7:0]    resultStage_controlPipeBeforePipe_s2mPipe_rData_horizontalDiff;
  reg        [7:0]    resultStage_controlPipeBeforePipe_s2mPipe_rData_verticalDiff;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_isHorizontalMin;
  reg        [7:0]    resultStage_controlPipeBeforePipe_s2mPipe_rData_minDiff;
  reg        [1:0]    resultStage_controlPipeBeforePipe_s2mPipe_rData_currentPosition;
  reg        [1:0]    resultStage_controlPipeBeforePipe_s2mPipe_rData_nextPosition;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_horizontalDirectionValid;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_verticalDirectionValid;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_mainDirectionValid;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_counterDirectionValid;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_inValidMinDiff;
  wire                when_Stream_l368_66;
  wire                resultStage_pixelStream_valid;
  wire                resultStage_pixelStream_ready;
  reg        [7:0]    resultStage_pixelStream_payload;
  wire                when_SuperResolutionPart3_l840;
  wire                when_SuperResolutionPart3_l846;
  wire                when_SuperResolutionPart3_l847;
  wire                when_SuperResolutionPart3_l850;
  wire                when_SuperResolutionPart3_l854;
  wire                when_SuperResolutionPart3_l855;
  wire                when_SuperResolutionPart3_l860;
  wire                when_SuperResolutionPart3_l861;
  wire                when_SuperResolutionPart3_l851;
  wire                when_SuperResolutionPart3_l841;
  wire                when_SuperResolutionPart3_l842;
  wire                when_SuperResolutionPart3_l869;
  wire                when_SuperResolutionPart3_l870;
  wire                when_SuperResolutionPart3_l871;
  wire                when_SuperResolutionPart3_l872;
  wire                when_SuperResolutionPart3_l875;
  wire                when_SuperResolutionPart3_l876;
  wire                when_SuperResolutionPart3_l885;
  wire                when_SuperResolutionPart3_l893;
  wire                when_SuperResolutionPart3_l884;
  wire                when_SuperResolutionPart3_l902;
  wire                when_SuperResolutionPart3_l903;
  wire                when_SuperResolutionPart3_l912;
  wire                when_SuperResolutionPart3_l920;
  wire                when_SuperResolutionPart3_l911;
  wire                when_SuperResolutionPart3_l874;
  wire                when_SuperResolutionPart3_l930;
  wire                when_SuperResolutionPart3_l931;
  wire                when_SuperResolutionPart3_l932;
  wire                when_SuperResolutionPart3_l941;
  wire                when_SuperResolutionPart3_l949;
  wire                when_SuperResolutionPart3_l940;
  wire                when_SuperResolutionPart3_l958;
  wire                when_SuperResolutionPart3_l959;
  wire                when_SuperResolutionPart3_l968;
  wire                when_SuperResolutionPart3_l976;
  wire                when_SuperResolutionPart3_l967;
  wire                when_SuperResolutionPart3_l986;
  wire                when_SuperResolutionPart3_l987;
  wire                when_SuperResolutionPart3_l988;
  wire                when_SuperResolutionPart3_l991;
  wire                when_SuperResolutionPart3_l992;
  wire                when_SuperResolutionPart3_l1001;
  wire                when_SuperResolutionPart3_l1009;
  wire                when_SuperResolutionPart3_l1000;
  wire                when_SuperResolutionPart3_l1019;
  wire                when_SuperResolutionPart3_l1020;
  wire                when_SuperResolutionPart3_l1021;
  wire                when_SuperResolutionPart3_l1024;
  wire                when_SuperResolutionPart3_l1025;
  wire                when_SuperResolutionPart3_l1034;
  wire                when_SuperResolutionPart3_l1042;
  wire                when_SuperResolutionPart3_l1033;
  wire                when_SuperResolutionPart3_l1052;
  wire                when_SuperResolutionPart3_l1053;
  wire                when_SuperResolutionPart3_l1062;
  wire                when_SuperResolutionPart3_l1070;
  wire                when_SuperResolutionPart3_l1061;
  wire                when_SuperResolutionPart3_l1079;
  wire                when_SuperResolutionPart3_l1080;
  wire                when_SuperResolutionPart3_l1083;
  wire                when_SuperResolutionPart3_l1084;
  wire                when_SuperResolutionPart3_l1093;
  wire                when_SuperResolutionPart3_l1101;
  wire                when_SuperResolutionPart3_l1092;
  wire                when_SuperResolutionPart3_l929;
  wire                when_SuperResolutionPart3_l985;
  wire                when_SuperResolutionPart3_l1018;
  wire                when_SuperResolutionPart3_l1051;
  wire                when_SuperResolutionPart3_l1078;
  wire                when_SuperResolutionPart3_l1082;
  wire                resultStage_pixelStream_s2mPipe_valid;
  reg                 resultStage_pixelStream_s2mPipe_ready;
  wire       [7:0]    resultStage_pixelStream_s2mPipe_payload;
  reg                 resultStage_pixelStream_rValid;
  reg        [7:0]    resultStage_pixelStream_rData;
  wire                resultStage_resultStream_valid;
  wire                resultStage_resultStream_ready;
  wire       [7:0]    resultStage_resultStream_payload;
  reg                 resultStage_pixelStream_s2mPipe_rValid;
  reg        [7:0]    resultStage_pixelStream_s2mPipe_rData;
  wire                when_Stream_l368_67;
  wire                when_SuperResolutionPart3_l1115;
  wire                diffStage_controlPipe_fire;
  wire                CICC1851_resultStage_mainOnePixelStream_ready;
  reg                 CICC1851_resultStage_mainOnePixelStream_ready_1;
  wire                CICC1851_resultStage_mainOnePixelStream_ready_2;
  wire                when_Stream_l438;
  reg                 resultsJoin_valid;
  wire                resultsJoin_ready;
  wire                pixelsStream_valid;
  wire                pixelsStream_ready;
  wire       [7:0]    pixelsStream_payload_pixel;
  wire                pixelsStream_payload_frameStart;
  wire                pixelsStream_payload_rowEnd;
  wire                pixelsStream_s2mPipe_valid;
  reg                 pixelsStream_s2mPipe_ready;
  wire       [7:0]    pixelsStream_s2mPipe_payload_pixel;
  wire                pixelsStream_s2mPipe_payload_frameStart;
  wire                pixelsStream_s2mPipe_payload_rowEnd;
  reg                 pixelsStream_rValid;
  reg        [7:0]    pixelsStream_rData_pixel;
  reg                 pixelsStream_rData_frameStart;
  reg                 pixelsStream_rData_rowEnd;
  wire                pixelsStream_s2mPipe_m2sPipe_valid;
  wire                pixelsStream_s2mPipe_m2sPipe_ready;
  wire       [7:0]    pixelsStream_s2mPipe_m2sPipe_payload_pixel;
  wire                pixelsStream_s2mPipe_m2sPipe_payload_frameStart;
  wire                pixelsStream_s2mPipe_m2sPipe_payload_rowEnd;
  reg                 pixelsStream_s2mPipe_rValid;
  reg        [7:0]    pixelsStream_s2mPipe_rData_pixel;
  reg                 pixelsStream_s2mPipe_rData_frameStart;
  reg                 pixelsStream_s2mPipe_rData_rowEnd;
  wire                when_Stream_l368_68;
  wire                controlStateMachine_wantExit;
  reg                 controlStateMachine_wantStart;
  wire                controlStateMachine_wantKill;
  reg        [1:0]    controlStateMachine_stateReg;
  reg        [1:0]    controlStateMachine_stateNext;
  wire                passPixels_fire_13;
  wire                when_SuperResolutionPart3_l1158;
  wire                controlStream_fire;
  wire                when_SuperResolutionPart3_l1168;
  wire                when_SuperResolutionPart3_l1188;
  wire                controlStream_fire_1;
  wire                when_SuperResolutionPart3_l1199;
  wire                passPixels_fire_14;
  wire                when_SuperResolutionPart3_l1202;
  wire                passPixels_fire_15;
  wire                when_SuperResolutionPart3_l1205;
  wire                when_SuperResolutionPart3_l1217;
  wire                controlStream_fire_2;
  wire                when_SuperResolutionPart3_l1220;
  wire                controlStream_fire_3;
  wire                when_SuperResolutionPart3_l1223;
  wire                controlStream_fire_4;
  wire                when_SuperResolutionPart3_l1224;
  wire                controlStream_fire_5;
  wire                when_SuperResolutionPart3_l1226;
  wire                controlStream_fire_6;
  wire                controlStream_fire_7;
  wire                when_SuperResolutionPart3_l1247;
  wire                when_SuperResolutionPart3_l1248;
  wire                when_SuperResolutionPart3_l1250;
  wire                when_SuperResolutionPart3_l1252;
  `ifndef SYNTHESIS
  reg [39:0] controlStateMachine_stateReg_string;
  reg [39:0] controlStateMachine_stateNext_string;
  `endif

  reg [7:0] lineBufferOne [0:3839];
  reg [7:0] lineBufferTwo [0:3839];
  reg [7:0] lineBufferThree [0:3839];
  reg [0:0] validBufferOne [0:3839];
  reg [0:0] validBufferTwo [0:3839];
  reg [0:0] validBufferThree [0:3839];

  assign CICC1851_bufferRowCount_valueNext_1 = bufferRowCount_willIncrement;
  assign CICC1851_bufferRowCount_valueNext = {11'd0, CICC1851_bufferRowCount_valueNext_1};
  assign CICC1851_bufferWAddr_valueNext_1 = bufferWAddr_willIncrement;
  assign CICC1851_bufferWAddr_valueNext = {11'd0, CICC1851_bufferWAddr_valueNext_1};
  assign CICC1851_outPixelAddr_valueNext_1 = outPixelAddr_willIncrement;
  assign CICC1851_outPixelAddr_valueNext = {11'd0, CICC1851_outPixelAddr_valueNext_1};
  assign CICC1851_outRowCount_valueNext_1 = outRowCount_willIncrement;
  assign CICC1851_outRowCount_valueNext = {11'd0, CICC1851_outRowCount_valueNext_1};
  assign CICC1851_alreadySendRow_valueNext_1 = alreadySendRow_willIncrement;
  assign CICC1851_alreadySendRow_valueNext = {11'd0, CICC1851_alreadySendRow_valueNext_1};
  assign CICC1851_alreadySendCountInRow_valueNext_1 = alreadySendCountInRow_willIncrement;
  assign CICC1851_alreadySendCountInRow_valueNext = {11'd0, CICC1851_alreadySendCountInRow_valueNext_1};
  assign CICC1851_nextRowBuffer = 1'b1;
  assign CICC1851_when_SuperResolutionPart3_l226 = {1'd0, bufferWAddr_value};
  assign CICC1851_when_SuperResolutionPart3_l226_1 = (CICC1851_when_SuperResolutionPart3_l226_2 - 13'h0002);
  assign CICC1851_when_SuperResolutionPart3_l226_2 = (3'b100 * bmpWidth);
  assign CICC1851_when_SuperResolutionPart3_l227 = {1'd0, bufferRowCount_value};
  assign CICC1851_when_SuperResolutionPart3_l227_1 = (CICC1851_when_SuperResolutionPart3_l227_2 - 13'h0002);
  assign CICC1851_when_SuperResolutionPart3_l227_2 = (3'b100 * bmpHeight);
  assign CICC1851_when_SuperResolutionPart3_l270 = {1'd0, alreadySendCountInRow_value};
  assign CICC1851_when_SuperResolutionPart3_l270_1 = (CICC1851_when_SuperResolutionPart3_l270_2 - 13'h0002);
  assign CICC1851_when_SuperResolutionPart3_l270_2 = (3'b100 * bmpWidth);
  assign CICC1851_when_SuperResolutionPart3_l271 = {1'd0, alreadySendRow_value};
  assign CICC1851_when_SuperResolutionPart3_l271_1 = (CICC1851_when_SuperResolutionPart3_l271_2 - 13'h0002);
  assign CICC1851_when_SuperResolutionPart3_l271_2 = (3'b100 * bmpHeight);
  assign CICC1851_resultStage_pixelStream_payload = (CICC1851_resultStage_pixelStream_payload_1 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_1 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_mainThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_2 = (CICC1851_resultStage_pixelStream_payload_3 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_3 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_mainThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_4 = (CICC1851_resultStage_pixelStream_payload_5 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_5 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_mainTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_6 = (CICC1851_resultStage_pixelStream_payload_7 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_7 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_mainThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_8 = (CICC1851_resultStage_pixelStream_payload_9 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_9 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_mainThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_10 = (CICC1851_resultStage_pixelStream_payload_11 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_11 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_mainTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_12 = (CICC1851_resultStage_pixelStream_payload_13 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_13 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_mainThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_14 = (CICC1851_resultStage_pixelStream_payload_15 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_15 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_mainThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_16 = (CICC1851_resultStage_pixelStream_payload_17 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_17 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_mainTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_18 = (CICC1851_resultStage_pixelStream_payload_19 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_19 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_20 = (CICC1851_resultStage_pixelStream_payload_21 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_21 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_22 = (CICC1851_resultStage_pixelStream_payload_23 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_23 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_24 = (CICC1851_resultStage_pixelStream_payload_25 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_25 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_26 = (CICC1851_resultStage_pixelStream_payload_27 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_27 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_28 = (CICC1851_resultStage_pixelStream_payload_29 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_29 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_30 = (CICC1851_resultStage_pixelStream_payload_31 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_31 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_32 = (CICC1851_resultStage_pixelStream_payload_33 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_33 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_34 = (CICC1851_resultStage_pixelStream_payload_35 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_35 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_36 = (CICC1851_resultStage_pixelStream_payload_37 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_37 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_38 = (CICC1851_resultStage_pixelStream_payload_39 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_39 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_40 = (CICC1851_resultStage_pixelStream_payload_41 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_41 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_42 = (CICC1851_resultStage_pixelStream_payload_43 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_43 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_44 = (CICC1851_resultStage_pixelStream_payload_45 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_45 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_46 = (CICC1851_resultStage_pixelStream_payload_47 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_47 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_48 = (CICC1851_resultStage_pixelStream_payload_49 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_49 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_50 = (CICC1851_resultStage_pixelStream_payload_51 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_51 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_52 = (CICC1851_resultStage_pixelStream_payload_53 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_53 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_54 = (CICC1851_resultStage_pixelStream_payload_55 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_55 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_56 = (CICC1851_resultStage_pixelStream_payload_57 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_57 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_58 = (CICC1851_resultStage_pixelStream_payload_59 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_59 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_60 = (CICC1851_resultStage_pixelStream_payload_61 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_61 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_62 = (CICC1851_resultStage_pixelStream_payload_63 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_63 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_64 = (CICC1851_resultStage_pixelStream_payload_65 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_65 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_66 = (CICC1851_resultStage_pixelStream_payload_67 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_67 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_68 = (CICC1851_resultStage_pixelStream_payload_69 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_69 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_70 = (CICC1851_resultStage_pixelStream_payload_71 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_71 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_72 = (CICC1851_resultStage_pixelStream_payload_73 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_73 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_74 = (CICC1851_resultStage_pixelStream_payload_75 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_75 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_76 = (CICC1851_resultStage_pixelStream_payload_77 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_77 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_78 = (CICC1851_resultStage_pixelStream_payload_79 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_79 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_80 = (CICC1851_resultStage_pixelStream_payload_81 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_81 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_82 = (CICC1851_resultStage_pixelStream_payload_83 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_83 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_84 = (CICC1851_resultStage_pixelStream_payload_85 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_85 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_86 = (CICC1851_resultStage_pixelStream_payload_87 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_87 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_88 = (CICC1851_resultStage_pixelStream_payload_89 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_89 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_90 = (CICC1851_resultStage_pixelStream_payload_91 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_91 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_92 = (CICC1851_resultStage_pixelStream_payload_93 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_93 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_94 = (CICC1851_resultStage_pixelStream_payload_95 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_95 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_96 = (CICC1851_resultStage_pixelStream_payload_97 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_97 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_98 = (CICC1851_resultStage_pixelStream_payload_99 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_99 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_100 = (CICC1851_resultStage_pixelStream_payload_101 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_101 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_102 = (CICC1851_resultStage_pixelStream_payload_103 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_103 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_104 = (CICC1851_resultStage_pixelStream_payload_105 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_105 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_106 = (CICC1851_resultStage_pixelStream_payload_107 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_107 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_108 = (CICC1851_resultStage_pixelStream_payload_109 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_109 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_110 = (CICC1851_resultStage_pixelStream_payload_111 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_111 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_112 = (CICC1851_resultStage_pixelStream_payload_113 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_113 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_114 = (CICC1851_resultStage_pixelStream_payload_115 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_115 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_116 = (CICC1851_resultStage_pixelStream_payload_117 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_117 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_118 = (CICC1851_resultStage_pixelStream_payload_119 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_119 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_120 = (CICC1851_resultStage_pixelStream_payload_121 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_121 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_122 = (CICC1851_resultStage_pixelStream_payload_123 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_123 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_124 = (CICC1851_resultStage_pixelStream_payload_125 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_125 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_126 = (CICC1851_resultStage_pixelStream_payload_127 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_127 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_128 = (CICC1851_resultStage_pixelStream_payload_129 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_129 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_130 = (CICC1851_resultStage_pixelStream_payload_131 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_131 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_132 = (CICC1851_resultStage_pixelStream_payload_133 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_133 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_134 = (CICC1851_resultStage_pixelStream_payload_135 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_135 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_136 = (CICC1851_resultStage_pixelStream_payload_137 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_137 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_138 = (CICC1851_resultStage_pixelStream_payload_139 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_139 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_140 = (CICC1851_resultStage_pixelStream_payload_141 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_141 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_142 = (CICC1851_resultStage_pixelStream_payload_143 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_143 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_144 = (CICC1851_resultStage_pixelStream_payload_145 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_145 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_146 = (CICC1851_resultStage_pixelStream_payload_147 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_147 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_148 = (CICC1851_resultStage_pixelStream_payload_149 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_149 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_150 = (CICC1851_resultStage_pixelStream_payload_151 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_151 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_152 = (CICC1851_resultStage_pixelStream_payload_153 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_153 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_154 = (CICC1851_resultStage_pixelStream_payload_155 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_155 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_156 = (CICC1851_resultStage_pixelStream_payload_157 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_157 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_158 = (CICC1851_resultStage_pixelStream_payload_159 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_159 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_160 = (CICC1851_resultStage_pixelStream_payload_161 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_161 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_162 = (CICC1851_resultStage_pixelStream_payload_163 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_163 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_164 = (CICC1851_resultStage_pixelStream_payload_165 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_165 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_166 = (CICC1851_resultStage_pixelStream_payload_167 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_167 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_168 = (CICC1851_resultStage_pixelStream_payload_169 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_169 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_170 = (CICC1851_resultStage_pixelStream_payload_171 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_171 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_172 = (CICC1851_resultStage_pixelStream_payload_173 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_173 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_174 = (CICC1851_resultStage_pixelStream_payload_175 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_175 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_176 = (CICC1851_resultStage_pixelStream_payload_177 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_177 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_178 = (CICC1851_resultStage_pixelStream_payload_179 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_179 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_180 = (CICC1851_resultStage_pixelStream_payload_181 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_181 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_182 = (CICC1851_resultStage_pixelStream_payload_183 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_183 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_184 = (CICC1851_resultStage_pixelStream_payload_185 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_185 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_186 = (CICC1851_resultStage_pixelStream_payload_187 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_187 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_188 = (CICC1851_resultStage_pixelStream_payload_189 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_189 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_190 = (CICC1851_resultStage_pixelStream_payload_191 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_191 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_192 = (CICC1851_resultStage_pixelStream_payload_193 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_193 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_194 = (CICC1851_resultStage_pixelStream_payload_195 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_195 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_196 = (CICC1851_resultStage_pixelStream_payload_197 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_197 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_198 = (CICC1851_resultStage_pixelStream_payload_199 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_199 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_200 = (CICC1851_resultStage_pixelStream_payload_201 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_201 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_202 = (CICC1851_resultStage_pixelStream_payload_203 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_203 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_204 = (CICC1851_resultStage_pixelStream_payload_205 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_205 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_206 = (CICC1851_resultStage_pixelStream_payload_207 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_207 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_208 = (CICC1851_resultStage_pixelStream_payload_209 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_209 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_210 = (CICC1851_resultStage_pixelStream_payload_211 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_211 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_212 = (CICC1851_resultStage_pixelStream_payload_213 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_213 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_214 = (CICC1851_resultStage_pixelStream_payload_215 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_215 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_216 = (CICC1851_resultStage_pixelStream_payload_217 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_217 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_218 = (CICC1851_resultStage_pixelStream_payload_219 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_219 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_220 = (CICC1851_resultStage_pixelStream_payload_221 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_221 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_222 = (CICC1851_resultStage_pixelStream_payload_223 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_223 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_224 = (CICC1851_resultStage_pixelStream_payload_225 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_225 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_226 = (CICC1851_resultStage_pixelStream_payload_227 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_227 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_228 = (CICC1851_resultStage_pixelStream_payload_229 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_229 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_230 = (CICC1851_resultStage_pixelStream_payload_231 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_231 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_232 = (CICC1851_resultStage_pixelStream_payload_233 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_233 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_234 = (CICC1851_resultStage_pixelStream_payload_235 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_235 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_236 = (CICC1851_resultStage_pixelStream_payload_237 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_237 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_238 = (CICC1851_resultStage_pixelStream_payload_239 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_239 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_240 = (CICC1851_resultStage_pixelStream_payload_241 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_241 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_242 = (CICC1851_resultStage_pixelStream_payload_243 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_243 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_244 = (CICC1851_resultStage_pixelStream_payload_245 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_245 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_246 = (CICC1851_resultStage_pixelStream_payload_247 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_247 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_248 = (CICC1851_resultStage_pixelStream_payload_249 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_249 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_when_SuperResolutionPart3_l1202 = (12'h003 + outRowCount_value);
  assign CICC1851_when_SuperResolutionPart3_l1205 = (12'h001 + outRowCount_value);
  assign CICC1851_when_SuperResolutionPart3_l1205_1 = (12'h002 + outPixelAddr_value);
  assign CICC1851_when_SuperResolutionPart3_l1205_2 = (12'h002 + outPixelAddr_value);
  assign CICC1851_when_SuperResolutionPart3_l1223 = {1'd0, outPixelAddr_value};
  assign CICC1851_when_SuperResolutionPart3_l1223_1 = (CICC1851_when_SuperResolutionPart3_l1223_2 - 13'h0002);
  assign CICC1851_when_SuperResolutionPart3_l1223_2 = (3'b100 * bmpWidth);
  assign CICC1851_when_SuperResolutionPart3_l1224 = {1'd0, outRowCount_value};
  assign CICC1851_when_SuperResolutionPart3_l1224_1 = (CICC1851_when_SuperResolutionPart3_l1224_2 - 13'h0002);
  assign CICC1851_when_SuperResolutionPart3_l1224_2 = (3'b100 * bmpHeight);
  assign CICC1851_lineBufferOne_port = passPixels_payload_pixel;
  assign CICC1851_lineBufferOne_port_1 = (passPixels_fire_6 && (bufferSwitch == 2'b00));
  assign CICC1851_lineBufferTwo_port = passPixels_payload_pixel;
  assign CICC1851_lineBufferTwo_port_1 = (passPixels_fire_7 && (bufferSwitch == 2'b01));
  assign CICC1851_lineBufferThree_port = passPixels_payload_pixel;
  assign CICC1851_lineBufferThree_port_1 = (passPixels_fire_8 && (bufferSwitch == 2'b10));
  assign CICC1851_validBufferOne_port = passPixels_payload_inpValid;
  assign CICC1851_validBufferOne_port_1 = (passPixels_fire_9 && (bufferSwitch == 2'b00));
  assign CICC1851_validBufferTwo_port = passPixels_payload_inpValid;
  assign CICC1851_validBufferTwo_port_1 = (passPixels_fire_10 && (bufferSwitch == 2'b01));
  assign CICC1851_validBufferThree_port = passPixels_payload_inpValid;
  assign CICC1851_validBufferThree_port_1 = (passPixels_fire_11 && (bufferSwitch == 2'b10));
  always @(posedge clk) begin
    if(CICC1851_lineBufferOne_port_1) begin
      lineBufferOne[bufferWAddr_value] <= CICC1851_lineBufferOne_port;
    end
  end

  always @(posedge clk) begin
    if(mainPixelAddrOneStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferOne_port1 <= lineBufferOne[mainPixelAddrOneStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(counterPixelAddrOneStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferOne_port2 <= lineBufferOne[counterPixelAddrOneStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(CICC1851_lineBufferTwo_port_1) begin
      lineBufferTwo[bufferWAddr_value] <= CICC1851_lineBufferTwo_port;
    end
  end

  always @(posedge clk) begin
    if(mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferTwo_port1 <= lineBufferTwo[mainPixelAddrTwoStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferTwo_port2 <= lineBufferTwo[counterPixelAddrTwoStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(CICC1851_lineBufferThree_port_1) begin
      lineBufferThree[bufferWAddr_value] <= CICC1851_lineBufferThree_port;
    end
  end

  always @(posedge clk) begin
    if(mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferThree_port1 <= lineBufferThree[mainPixelAddrThreeStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferThree_port2 <= lineBufferThree[counterPixelAddrThreeStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(CICC1851_validBufferOne_port_1) begin
      validBufferOne[bufferWAddr_value] <= CICC1851_validBufferOne_port;
    end
  end

  always @(posedge clk) begin
    if(mainValidAddrOneStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_validBufferOne_port1 <= validBufferOne[mainValidAddrOneStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(counterValidAddrOneStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_validBufferOne_port2 <= validBufferOne[counterValidAddrOneStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(CICC1851_validBufferTwo_port_1) begin
      validBufferTwo[bufferWAddr_value] <= CICC1851_validBufferTwo_port;
    end
  end

  always @(posedge clk) begin
    if(mainValidAddrTwoStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_validBufferTwo_port1 <= validBufferTwo[mainValidAddrTwoStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(counterValidAddrTwoStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_validBufferTwo_port2 <= validBufferTwo[counterValidAddrTwoStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(CICC1851_validBufferThree_port_1) begin
      validBufferThree[bufferWAddr_value] <= CICC1851_validBufferThree_port;
    end
  end

  always @(posedge clk) begin
    if(mainValidAddrThreeStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_validBufferThree_port1 <= validBufferThree[mainValidAddrThreeStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(counterValidAddrThreeStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_validBufferThree_port2 <= validBufferThree[counterValidAddrThreeStream_s2mPipe_m2sPipe_payload];
    end
  end

  StreamFork_3 diffStage_controlPipe_fork (
    .io_input_valid                                (diffStage_controlPipe_valid                                             ), //i
    .io_input_ready                                (diffStage_controlPipe_fork_io_input_ready                               ), //o
    .io_input_payload_frameStart                   (diffStage_controlPipe_payload_frameStart                                ), //i
    .io_input_payload_rowEnd                       (diffStage_controlPipe_payload_rowEnd                                    ), //i
    .io_input_payload_pipeValid                    (diffStage_controlPipe_payload_pipeValid                                 ), //i
    .io_input_payload_firstRow                     (diffStage_controlPipe_payload_firstRow                                  ), //i
    .io_input_payload_lastRow                      (diffStage_controlPipe_payload_lastRow                                   ), //i
    .io_input_payload_finalResult                  (diffStage_controlPipe_payload_finalResult                               ), //i
    .io_input_payload_mainCompare                  (diffStage_controlPipe_payload_mainCompare                               ), //i
    .io_input_payload_counterCompare               (diffStage_controlPipe_payload_counterCompare                            ), //i
    .io_input_payload_horizontalCompare            (diffStage_controlPipe_payload_horizontalCompare                         ), //i
    .io_input_payload_verticalCompare              (diffStage_controlPipe_payload_verticalCompare                           ), //i
    .io_input_payload_mainDiff                     (diffStage_controlPipe_payload_mainDiff[7:0]                             ), //i
    .io_input_payload_counterDiff                  (diffStage_controlPipe_payload_counterDiff[7:0]                          ), //i
    .io_input_payload_horizontalDiff               (diffStage_controlPipe_payload_horizontalDiff[7:0]                       ), //i
    .io_input_payload_verticalDiff                 (diffStage_controlPipe_payload_verticalDiff[7:0]                         ), //i
    .io_input_payload_isHorizontalMin              (diffStage_controlPipe_payload_isHorizontalMin                           ), //i
    .io_input_payload_minDiff                      (diffStage_controlPipe_payload_minDiff[7:0]                              ), //i
    .io_input_payload_currentPosition              (diffStage_controlPipe_payload_currentPosition[1:0]                      ), //i
    .io_input_payload_nextPosition                 (diffStage_controlPipe_payload_nextPosition[1:0]                         ), //i
    .io_input_payload_horizontalDirectionValid     (diffStage_controlPipe_payload_horizontalDirectionValid                  ), //i
    .io_input_payload_verticalDirectionValid       (diffStage_controlPipe_payload_verticalDirectionValid                    ), //i
    .io_input_payload_mainDirectionValid           (diffStage_controlPipe_payload_mainDirectionValid                        ), //i
    .io_input_payload_counterDirectionValid        (diffStage_controlPipe_payload_counterDirectionValid                     ), //i
    .io_input_payload_inValidMinDiff               (diffStage_controlPipe_payload_inValidMinDiff                            ), //i
    .io_outputs_0_valid                            (diffStage_controlPipe_fork_io_outputs_0_valid                           ), //o
    .io_outputs_0_ready                            (resultStage_controlPipeBeforePipe_ready                                 ), //i
    .io_outputs_0_payload_frameStart               (diffStage_controlPipe_fork_io_outputs_0_payload_frameStart              ), //o
    .io_outputs_0_payload_rowEnd                   (diffStage_controlPipe_fork_io_outputs_0_payload_rowEnd                  ), //o
    .io_outputs_0_payload_pipeValid                (diffStage_controlPipe_fork_io_outputs_0_payload_pipeValid               ), //o
    .io_outputs_0_payload_firstRow                 (diffStage_controlPipe_fork_io_outputs_0_payload_firstRow                ), //o
    .io_outputs_0_payload_lastRow                  (diffStage_controlPipe_fork_io_outputs_0_payload_lastRow                 ), //o
    .io_outputs_0_payload_finalResult              (diffStage_controlPipe_fork_io_outputs_0_payload_finalResult             ), //o
    .io_outputs_0_payload_mainCompare              (diffStage_controlPipe_fork_io_outputs_0_payload_mainCompare             ), //o
    .io_outputs_0_payload_counterCompare           (diffStage_controlPipe_fork_io_outputs_0_payload_counterCompare          ), //o
    .io_outputs_0_payload_horizontalCompare        (diffStage_controlPipe_fork_io_outputs_0_payload_horizontalCompare       ), //o
    .io_outputs_0_payload_verticalCompare          (diffStage_controlPipe_fork_io_outputs_0_payload_verticalCompare         ), //o
    .io_outputs_0_payload_mainDiff                 (diffStage_controlPipe_fork_io_outputs_0_payload_mainDiff[7:0]           ), //o
    .io_outputs_0_payload_counterDiff              (diffStage_controlPipe_fork_io_outputs_0_payload_counterDiff[7:0]        ), //o
    .io_outputs_0_payload_horizontalDiff           (diffStage_controlPipe_fork_io_outputs_0_payload_horizontalDiff[7:0]     ), //o
    .io_outputs_0_payload_verticalDiff             (diffStage_controlPipe_fork_io_outputs_0_payload_verticalDiff[7:0]       ), //o
    .io_outputs_0_payload_isHorizontalMin          (diffStage_controlPipe_fork_io_outputs_0_payload_isHorizontalMin         ), //o
    .io_outputs_0_payload_minDiff                  (diffStage_controlPipe_fork_io_outputs_0_payload_minDiff[7:0]            ), //o
    .io_outputs_0_payload_currentPosition          (diffStage_controlPipe_fork_io_outputs_0_payload_currentPosition[1:0]    ), //o
    .io_outputs_0_payload_nextPosition             (diffStage_controlPipe_fork_io_outputs_0_payload_nextPosition[1:0]       ), //o
    .io_outputs_0_payload_horizontalDirectionValid (diffStage_controlPipe_fork_io_outputs_0_payload_horizontalDirectionValid), //o
    .io_outputs_0_payload_verticalDirectionValid   (diffStage_controlPipe_fork_io_outputs_0_payload_verticalDirectionValid  ), //o
    .io_outputs_0_payload_mainDirectionValid       (diffStage_controlPipe_fork_io_outputs_0_payload_mainDirectionValid      ), //o
    .io_outputs_0_payload_counterDirectionValid    (diffStage_controlPipe_fork_io_outputs_0_payload_counterDirectionValid   ), //o
    .io_outputs_0_payload_inValidMinDiff           (diffStage_controlPipe_fork_io_outputs_0_payload_inValidMinDiff          ), //o
    .io_outputs_1_valid                            (diffStage_controlPipe_fork_io_outputs_1_valid                           ), //o
    .io_outputs_1_ready                            (resultStage_pixelStream_ready                                           ), //i
    .io_outputs_1_payload_frameStart               (diffStage_controlPipe_fork_io_outputs_1_payload_frameStart              ), //o
    .io_outputs_1_payload_rowEnd                   (diffStage_controlPipe_fork_io_outputs_1_payload_rowEnd                  ), //o
    .io_outputs_1_payload_pipeValid                (diffStage_controlPipe_fork_io_outputs_1_payload_pipeValid               ), //o
    .io_outputs_1_payload_firstRow                 (diffStage_controlPipe_fork_io_outputs_1_payload_firstRow                ), //o
    .io_outputs_1_payload_lastRow                  (diffStage_controlPipe_fork_io_outputs_1_payload_lastRow                 ), //o
    .io_outputs_1_payload_finalResult              (diffStage_controlPipe_fork_io_outputs_1_payload_finalResult             ), //o
    .io_outputs_1_payload_mainCompare              (diffStage_controlPipe_fork_io_outputs_1_payload_mainCompare             ), //o
    .io_outputs_1_payload_counterCompare           (diffStage_controlPipe_fork_io_outputs_1_payload_counterCompare          ), //o
    .io_outputs_1_payload_horizontalCompare        (diffStage_controlPipe_fork_io_outputs_1_payload_horizontalCompare       ), //o
    .io_outputs_1_payload_verticalCompare          (diffStage_controlPipe_fork_io_outputs_1_payload_verticalCompare         ), //o
    .io_outputs_1_payload_mainDiff                 (diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff[7:0]           ), //o
    .io_outputs_1_payload_counterDiff              (diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff[7:0]        ), //o
    .io_outputs_1_payload_horizontalDiff           (diffStage_controlPipe_fork_io_outputs_1_payload_horizontalDiff[7:0]     ), //o
    .io_outputs_1_payload_verticalDiff             (diffStage_controlPipe_fork_io_outputs_1_payload_verticalDiff[7:0]       ), //o
    .io_outputs_1_payload_isHorizontalMin          (diffStage_controlPipe_fork_io_outputs_1_payload_isHorizontalMin         ), //o
    .io_outputs_1_payload_minDiff                  (diffStage_controlPipe_fork_io_outputs_1_payload_minDiff[7:0]            ), //o
    .io_outputs_1_payload_currentPosition          (diffStage_controlPipe_fork_io_outputs_1_payload_currentPosition[1:0]    ), //o
    .io_outputs_1_payload_nextPosition             (diffStage_controlPipe_fork_io_outputs_1_payload_nextPosition[1:0]       ), //o
    .io_outputs_1_payload_horizontalDirectionValid (diffStage_controlPipe_fork_io_outputs_1_payload_horizontalDirectionValid), //o
    .io_outputs_1_payload_verticalDirectionValid   (diffStage_controlPipe_fork_io_outputs_1_payload_verticalDirectionValid  ), //o
    .io_outputs_1_payload_mainDirectionValid       (diffStage_controlPipe_fork_io_outputs_1_payload_mainDirectionValid      ), //o
    .io_outputs_1_payload_counterDirectionValid    (diffStage_controlPipe_fork_io_outputs_1_payload_counterDirectionValid   ), //o
    .io_outputs_1_payload_inValidMinDiff           (diffStage_controlPipe_fork_io_outputs_1_payload_inValidMinDiff          )  //o
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_5_BOOT : controlStateMachine_stateReg_string = "BOOT ";
      controlStateMachine_enumDef_5_HOLD : controlStateMachine_stateReg_string = "HOLD ";
      controlStateMachine_enumDef_5_PASS : controlStateMachine_stateReg_string = "PASS ";
      controlStateMachine_enumDef_5_EXTRA : controlStateMachine_stateReg_string = "EXTRA";
      default : controlStateMachine_stateReg_string = "?????";
    endcase
  end
  always @(*) begin
    case(controlStateMachine_stateNext)
      controlStateMachine_enumDef_5_BOOT : controlStateMachine_stateNext_string = "BOOT ";
      controlStateMachine_enumDef_5_HOLD : controlStateMachine_stateNext_string = "HOLD ";
      controlStateMachine_enumDef_5_PASS : controlStateMachine_stateNext_string = "PASS ";
      controlStateMachine_enumDef_5_EXTRA : controlStateMachine_stateNext_string = "EXTRA";
      default : controlStateMachine_stateNext_string = "?????";
    endcase
  end
  `endif

  always @(*) begin
    pixelsIn_ready = 1'b0;
    pixelsIn_ready = (! pixelsIn_rValid);
  end

  always @(*) begin
    pixelsOut_valid = 1'b0;
    pixelsOut_valid = pixelsStream_s2mPipe_m2sPipe_valid;
  end

  always @(*) begin
    pixelsOut_payload_pixel = 8'h0;
    pixelsOut_payload_pixel = pixelsStream_s2mPipe_m2sPipe_payload_pixel;
  end

  always @(*) begin
    pixelsOut_payload_frameStart = 1'b0;
    pixelsOut_payload_frameStart = pixelsStream_s2mPipe_m2sPipe_payload_frameStart;
  end

  always @(*) begin
    pixelsOut_payload_rowEnd = 1'b0;
    pixelsOut_payload_rowEnd = pixelsStream_s2mPipe_m2sPipe_payload_rowEnd;
  end

  always @(*) begin
    inpThreeDoneOut = 1'b0;
    inpThreeDoneOut = inpThreeDone;
  end

  assign when_SuperResolutionPart3_l72 = (startIn && (! startIn_regNext));
  assign when_SuperResolutionPart3_l75 = (! startIn);
  assign when_SuperResolutionPart3_l78 = (startIn && (! readDone));
  assign when_SuperResolutionPart3_l78_1 = (! startIn);
  assign when_SuperResolutionPart3_l93 = (! startIn);
  assign when_SuperResolutionPart3_l96 = (! startIn);
  always @(*) begin
    bufferRowCount_willIncrement = 1'b0;
    if(when_SuperResolutionPart3_l230) begin
      if(!bufferReachFinalRow) begin
        bufferRowCount_willIncrement = 1'b1;
      end
    end
  end

  always @(*) begin
    bufferRowCount_willClear = 1'b0;
    if(when_SuperResolutionPart3_l230) begin
      if(bufferReachFinalRow) begin
        bufferRowCount_willClear = 1'b1;
      end
    end
  end

  assign bufferRowCount_willOverflowIfInc = (bufferRowCount_value == 12'h870);
  assign bufferRowCount_willOverflow = (bufferRowCount_willOverflowIfInc && bufferRowCount_willIncrement);
  always @(*) begin
    if(bufferRowCount_willOverflow) begin
      bufferRowCount_valueNext = 12'h0;
    end else begin
      bufferRowCount_valueNext = (bufferRowCount_value + CICC1851_bufferRowCount_valueNext);
    end
    if(bufferRowCount_willClear) begin
      bufferRowCount_valueNext = 12'h0;
    end
  end

  assign when_SuperResolutionPart3_l102 = ((startIn && (! holdBuffer)) && (! writeDone));
  assign when_SuperResolutionPart3_l102_1 = (((! startIn) || holdBuffer) || writeDone);
  always @(*) begin
    bufferWAddr_willIncrement = 1'b0;
    if(passPixels_fire_12) begin
      if(!passPixels_payload_rowEnd) begin
        bufferWAddr_willIncrement = 1'b1;
      end
    end
  end

  always @(*) begin
    bufferWAddr_willClear = 1'b0;
    if(passPixels_fire_12) begin
      if(passPixels_payload_rowEnd) begin
        bufferWAddr_willClear = 1'b1;
      end
    end
  end

  assign bufferWAddr_willOverflowIfInc = (bufferWAddr_value == 12'heff);
  assign bufferWAddr_willOverflow = (bufferWAddr_willOverflowIfInc && bufferWAddr_willIncrement);
  always @(*) begin
    if(bufferWAddr_willOverflow) begin
      bufferWAddr_valueNext = 12'h0;
    end else begin
      bufferWAddr_valueNext = (bufferWAddr_value + CICC1851_bufferWAddr_valueNext);
    end
    if(bufferWAddr_willClear) begin
      bufferWAddr_valueNext = 12'h0;
    end
  end

  always @(*) begin
    outPixelAddr_willIncrement = 1'b0;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_5_HOLD : begin
      end
      controlStateMachine_enumDef_5_PASS : begin
      end
      controlStateMachine_enumDef_5_EXTRA : begin
        if(controlStream_fire_6) begin
          if(!outReachRowEnd) begin
            outPixelAddr_willIncrement = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outPixelAddr_willClear = 1'b0;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_5_HOLD : begin
      end
      controlStateMachine_enumDef_5_PASS : begin
      end
      controlStateMachine_enumDef_5_EXTRA : begin
        if(controlStream_fire_6) begin
          if(outReachRowEnd) begin
            outPixelAddr_willClear = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign outPixelAddr_willOverflowIfInc = (outPixelAddr_value == 12'heff);
  assign outPixelAddr_willOverflow = (outPixelAddr_willOverflowIfInc && outPixelAddr_willIncrement);
  always @(*) begin
    if(outPixelAddr_willOverflow) begin
      outPixelAddr_valueNext = 12'h0;
    end else begin
      outPixelAddr_valueNext = (outPixelAddr_value + CICC1851_outPixelAddr_valueNext);
    end
    if(outPixelAddr_willClear) begin
      outPixelAddr_valueNext = 12'h0;
    end
  end

  always @(*) begin
    outRowCount_willIncrement = 1'b0;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_5_HOLD : begin
      end
      controlStateMachine_enumDef_5_PASS : begin
      end
      controlStateMachine_enumDef_5_EXTRA : begin
        if(when_SuperResolutionPart3_l1226) begin
          if(!outReachFinalRow) begin
            outRowCount_willIncrement = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outRowCount_willClear = 1'b0;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_5_HOLD : begin
      end
      controlStateMachine_enumDef_5_PASS : begin
      end
      controlStateMachine_enumDef_5_EXTRA : begin
        if(when_SuperResolutionPart3_l1226) begin
          if(outReachFinalRow) begin
            outRowCount_willClear = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign outRowCount_willOverflowIfInc = (outRowCount_value == 12'h870);
  assign outRowCount_willOverflow = (outRowCount_willOverflowIfInc && outRowCount_willIncrement);
  always @(*) begin
    if(outRowCount_willOverflow) begin
      outRowCount_valueNext = 12'h0;
    end else begin
      outRowCount_valueNext = (outRowCount_value + CICC1851_outRowCount_valueNext);
    end
    if(outRowCount_willClear) begin
      outRowCount_valueNext = 12'h0;
    end
  end

  always @(*) begin
    alreadySendRow_willIncrement = 1'b0;
    if(pixelsOut_fire_2) begin
      if(alreadyReachRowEnd) begin
        if(!alreadyReachFinalRow) begin
          alreadySendRow_willIncrement = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    alreadySendRow_willClear = 1'b0;
    if(pixelsOut_fire_2) begin
      if(alreadyReachRowEnd) begin
        if(alreadyReachFinalRow) begin
          alreadySendRow_willClear = 1'b1;
        end
      end
    end
  end

  assign alreadySendRow_willOverflowIfInc = (alreadySendRow_value == 12'h870);
  assign alreadySendRow_willOverflow = (alreadySendRow_willOverflowIfInc && alreadySendRow_willIncrement);
  always @(*) begin
    if(alreadySendRow_willOverflow) begin
      alreadySendRow_valueNext = 12'h0;
    end else begin
      alreadySendRow_valueNext = (alreadySendRow_value + CICC1851_alreadySendRow_valueNext);
    end
    if(alreadySendRow_willClear) begin
      alreadySendRow_valueNext = 12'h0;
    end
  end

  always @(*) begin
    alreadySendCountInRow_willIncrement = 1'b0;
    if(pixelsOut_fire_2) begin
      if(!alreadyReachRowEnd) begin
        alreadySendCountInRow_willIncrement = 1'b1;
      end
    end
  end

  always @(*) begin
    alreadySendCountInRow_willClear = 1'b0;
    if(pixelsOut_fire_2) begin
      if(alreadyReachRowEnd) begin
        alreadySendCountInRow_willClear = 1'b1;
      end
    end
  end

  assign alreadySendCountInRow_willOverflowIfInc = (alreadySendCountInRow_value == 12'heff);
  assign alreadySendCountInRow_willOverflow = (alreadySendCountInRow_willOverflowIfInc && alreadySendCountInRow_willIncrement);
  always @(*) begin
    if(alreadySendCountInRow_willOverflow) begin
      alreadySendCountInRow_valueNext = 12'h0;
    end else begin
      alreadySendCountInRow_valueNext = (alreadySendCountInRow_value + CICC1851_alreadySendCountInRow_valueNext);
    end
    if(alreadySendCountInRow_willClear) begin
      alreadySendCountInRow_valueNext = 12'h0;
    end
  end

  assign when_SuperResolutionPart3_l154 = ((! startRead) || ((! startIn) && startIn_regNext_1));
  always @(*) begin
    mainAddrOne = outPixelAddr_value;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_5_HOLD : begin
      end
      controlStateMachine_enumDef_5_PASS : begin
        if(when_SuperResolutionPart3_l1168) begin
          mainAddrOne = (12'h001 + outPixelAddr_value);
        end else begin
          mainAddrOne = (outPixelAddr_value - 12'h001);
        end
      end
      controlStateMachine_enumDef_5_EXTRA : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    counterAddrOne = outPixelAddr_value;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_5_HOLD : begin
      end
      controlStateMachine_enumDef_5_PASS : begin
        if(outReachRowEnd) begin
          counterAddrOne = (outPixelAddr_value - 12'h001);
        end else begin
          counterAddrOne = (12'h001 + outPixelAddr_value);
        end
      end
      controlStateMachine_enumDef_5_EXTRA : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    mainAddrTwo = outPixelAddr_value;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_5_HOLD : begin
      end
      controlStateMachine_enumDef_5_PASS : begin
        if(when_SuperResolutionPart3_l1168) begin
          mainAddrTwo = (12'h001 + outPixelAddr_value);
        end else begin
          mainAddrTwo = (outPixelAddr_value - 12'h001);
        end
      end
      controlStateMachine_enumDef_5_EXTRA : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    counterAddrTwo = outPixelAddr_value;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_5_HOLD : begin
      end
      controlStateMachine_enumDef_5_PASS : begin
        if(outReachRowEnd) begin
          counterAddrTwo = (outPixelAddr_value - 12'h001);
        end else begin
          counterAddrTwo = (12'h001 + outPixelAddr_value);
        end
      end
      controlStateMachine_enumDef_5_EXTRA : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    mainAddrThree = outPixelAddr_value;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_5_HOLD : begin
      end
      controlStateMachine_enumDef_5_PASS : begin
        if(when_SuperResolutionPart3_l1168) begin
          mainAddrThree = (12'h001 + outPixelAddr_value);
        end else begin
          mainAddrThree = (outPixelAddr_value - 12'h001);
        end
      end
      controlStateMachine_enumDef_5_EXTRA : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    counterAddrThree = outPixelAddr_value;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_5_HOLD : begin
      end
      controlStateMachine_enumDef_5_PASS : begin
        if(outReachRowEnd) begin
          counterAddrThree = (outPixelAddr_value - 12'h001);
        end else begin
          counterAddrThree = (12'h001 + outPixelAddr_value);
        end
      end
      controlStateMachine_enumDef_5_EXTRA : begin
      end
      default : begin
      end
    endcase
  end

  assign validStream_valid = 1'b1;
  assign CICC1851_controls_frameStart = 60'h0;
  always @(*) begin
    controls_frameStart = CICC1851_controls_frameStart[0];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_5_HOLD : begin
      end
      controlStateMachine_enumDef_5_PASS : begin
        if(frameStart) begin
          controls_frameStart = 1'b1;
        end
      end
      controlStateMachine_enumDef_5_EXTRA : begin
        if(frameStart) begin
          controls_frameStart = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_rowEnd = CICC1851_controls_frameStart[1];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_5_HOLD : begin
      end
      controlStateMachine_enumDef_5_PASS : begin
        if(outReachRowEnd) begin
          controls_rowEnd = 1'b1;
        end
      end
      controlStateMachine_enumDef_5_EXTRA : begin
        if(outReachRowEnd) begin
          controls_rowEnd = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_pipeValid = CICC1851_controls_frameStart[2];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_5_HOLD : begin
      end
      controlStateMachine_enumDef_5_PASS : begin
        controls_pipeValid = 1'b1;
      end
      controlStateMachine_enumDef_5_EXTRA : begin
        controls_pipeValid = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_firstRow = CICC1851_controls_frameStart[3];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_5_HOLD : begin
      end
      controlStateMachine_enumDef_5_PASS : begin
        if(when_SuperResolutionPart3_l1188) begin
          controls_firstRow = 1'b1;
        end
      end
      controlStateMachine_enumDef_5_EXTRA : begin
        if(when_SuperResolutionPart3_l1217) begin
          controls_firstRow = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_lastRow = CICC1851_controls_frameStart[4];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_5_HOLD : begin
      end
      controlStateMachine_enumDef_5_PASS : begin
        if(outReachFinalRow) begin
          controls_lastRow = 1'b1;
        end
      end
      controlStateMachine_enumDef_5_EXTRA : begin
        if(outReachFinalRow) begin
          controls_lastRow = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_finalResult = CICC1851_controls_frameStart[5];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_5_HOLD : begin
      end
      controlStateMachine_enumDef_5_PASS : begin
      end
      controlStateMachine_enumDef_5_EXTRA : begin
        controls_finalResult = 1'b1;
      end
      default : begin
      end
    endcase
  end

  assign controls_mainCompare = CICC1851_controls_frameStart[6];
  assign controls_counterCompare = CICC1851_controls_frameStart[7];
  assign controls_horizontalCompare = CICC1851_controls_frameStart[8];
  assign controls_verticalCompare = CICC1851_controls_frameStart[9];
  assign controls_mainDiff = CICC1851_controls_frameStart[17 : 10];
  assign controls_counterDiff = CICC1851_controls_frameStart[25 : 18];
  assign controls_horizontalDiff = CICC1851_controls_frameStart[33 : 26];
  assign controls_verticalDiff = CICC1851_controls_frameStart[41 : 34];
  assign controls_isHorizontalMin = CICC1851_controls_frameStart[42];
  assign controls_minDiff = CICC1851_controls_frameStart[50 : 43];
  always @(*) begin
    controls_currentPosition = CICC1851_controls_frameStart[52 : 51];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_5_HOLD : begin
      end
      controlStateMachine_enumDef_5_PASS : begin
        controls_currentPosition = currentRowBuffer;
      end
      controlStateMachine_enumDef_5_EXTRA : begin
        controls_currentPosition = currentRowBuffer;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_nextPosition = CICC1851_controls_frameStart[54 : 53];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_5_HOLD : begin
      end
      controlStateMachine_enumDef_5_PASS : begin
        controls_nextPosition = nextRowBuffer;
      end
      controlStateMachine_enumDef_5_EXTRA : begin
        controls_nextPosition = nextRowBuffer;
      end
      default : begin
      end
    endcase
  end

  assign controls_horizontalDirectionValid = CICC1851_controls_frameStart[55];
  assign controls_verticalDirectionValid = CICC1851_controls_frameStart[56];
  assign controls_mainDirectionValid = CICC1851_controls_frameStart[57];
  assign controls_counterDirectionValid = CICC1851_controls_frameStart[58];
  assign controls_inValidMinDiff = CICC1851_controls_frameStart[59];
  always @(*) begin
    validStream_ready = (controlStream_ready && startRead);
    validStream_ready = (mainPixelAddrOneStream_ready && startRead);
    validStream_ready = (counterPixelAddrOneStream_ready && startRead);
    validStream_ready = (mainPixelAddrTwoStream_ready && startRead);
    validStream_ready = (counterPixelAddrTwoStream_ready && startRead);
    validStream_ready = (mainPixelAddrThreeStream_ready && startRead);
    validStream_ready = (counterPixelAddrThreeStream_ready && startRead);
    validStream_ready = (mainValidAddrOneStream_ready && startRead);
    validStream_ready = (counterValidAddrOneStream_ready && startRead);
    validStream_ready = (mainValidAddrTwoStream_ready && startRead);
    validStream_ready = (counterValidAddrTwoStream_ready && startRead);
    validStream_ready = (mainValidAddrThreeStream_ready && startRead);
    validStream_ready = (counterValidAddrThreeStream_ready && startRead);
  end

  assign controlStream_valid = (validStream_valid && startRead);
  assign controlStream_payload_frameStart = controls_frameStart;
  assign controlStream_payload_rowEnd = controls_rowEnd;
  assign controlStream_payload_pipeValid = controls_pipeValid;
  assign controlStream_payload_firstRow = controls_firstRow;
  assign controlStream_payload_lastRow = controls_lastRow;
  assign controlStream_payload_finalResult = controls_finalResult;
  assign controlStream_payload_mainCompare = controls_mainCompare;
  assign controlStream_payload_counterCompare = controls_counterCompare;
  assign controlStream_payload_horizontalCompare = controls_horizontalCompare;
  assign controlStream_payload_verticalCompare = controls_verticalCompare;
  assign controlStream_payload_mainDiff = controls_mainDiff;
  assign controlStream_payload_counterDiff = controls_counterDiff;
  assign controlStream_payload_horizontalDiff = controls_horizontalDiff;
  assign controlStream_payload_verticalDiff = controls_verticalDiff;
  assign controlStream_payload_isHorizontalMin = controls_isHorizontalMin;
  assign controlStream_payload_minDiff = controls_minDiff;
  assign controlStream_payload_currentPosition = controls_currentPosition;
  assign controlStream_payload_nextPosition = controls_nextPosition;
  assign controlStream_payload_horizontalDirectionValid = controls_horizontalDirectionValid;
  assign controlStream_payload_verticalDirectionValid = controls_verticalDirectionValid;
  assign controlStream_payload_mainDirectionValid = controls_mainDirectionValid;
  assign controlStream_payload_counterDirectionValid = controls_counterDirectionValid;
  assign controlStream_payload_inValidMinDiff = controls_inValidMinDiff;
  assign mainPixelAddrOneStream_valid = (validStream_valid && startRead);
  assign mainPixelAddrOneStream_payload = mainAddrOne;
  assign counterPixelAddrOneStream_valid = (validStream_valid && startRead);
  assign counterPixelAddrOneStream_payload = counterAddrOne;
  assign mainPixelAddrTwoStream_valid = (validStream_valid && startRead);
  assign mainPixelAddrTwoStream_payload = mainAddrTwo;
  assign counterPixelAddrTwoStream_valid = (validStream_valid && startRead);
  assign counterPixelAddrTwoStream_payload = counterAddrTwo;
  assign mainPixelAddrThreeStream_valid = (validStream_valid && startRead);
  assign mainPixelAddrThreeStream_payload = mainAddrThree;
  assign counterPixelAddrThreeStream_valid = (validStream_valid && startRead);
  assign counterPixelAddrThreeStream_payload = counterAddrThree;
  assign mainValidAddrOneStream_valid = (validStream_valid && startRead);
  assign mainValidAddrOneStream_payload = mainAddrOne;
  assign counterValidAddrOneStream_valid = (validStream_valid && startRead);
  assign counterValidAddrOneStream_payload = counterAddrOne;
  assign mainValidAddrTwoStream_valid = (validStream_valid && startRead);
  assign mainValidAddrTwoStream_payload = mainAddrTwo;
  assign counterValidAddrTwoStream_valid = (validStream_valid && startRead);
  assign counterValidAddrTwoStream_payload = counterAddrTwo;
  assign mainValidAddrThreeStream_valid = (validStream_valid && startRead);
  assign mainValidAddrThreeStream_payload = mainAddrThree;
  assign counterValidAddrThreeStream_valid = (validStream_valid && startRead);
  assign counterValidAddrThreeStream_payload = counterAddrThree;
  assign pixelsIn_s2mPipe_valid = (pixelsIn_valid || pixelsIn_rValid);
  assign pixelsIn_s2mPipe_payload_pixel = (pixelsIn_rValid ? pixelsIn_rData_pixel : pixelsIn_payload_pixel);
  assign pixelsIn_s2mPipe_payload_frameStart = (pixelsIn_rValid ? pixelsIn_rData_frameStart : pixelsIn_payload_frameStart);
  assign pixelsIn_s2mPipe_payload_rowEnd = (pixelsIn_rValid ? pixelsIn_rData_rowEnd : pixelsIn_payload_rowEnd);
  assign pixelsIn_s2mPipe_payload_inpValid = (pixelsIn_rValid ? pixelsIn_rData_inpValid : pixelsIn_payload_inpValid);
  always @(*) begin
    pixelsIn_s2mPipe_ready = pixelsIn_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368) begin
      pixelsIn_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368 = (! pixelsIn_s2mPipe_m2sPipe_valid);
  assign pixelsIn_s2mPipe_m2sPipe_valid = pixelsIn_s2mPipe_rValid;
  assign pixelsIn_s2mPipe_m2sPipe_payload_pixel = pixelsIn_s2mPipe_rData_pixel;
  assign pixelsIn_s2mPipe_m2sPipe_payload_frameStart = pixelsIn_s2mPipe_rData_frameStart;
  assign pixelsIn_s2mPipe_m2sPipe_payload_rowEnd = pixelsIn_s2mPipe_rData_rowEnd;
  assign pixelsIn_s2mPipe_m2sPipe_payload_inpValid = pixelsIn_s2mPipe_rData_inpValid;
  assign passPixels_valid = (pixelsIn_s2mPipe_m2sPipe_valid && bufferEnable);
  assign pixelsIn_s2mPipe_m2sPipe_ready = (passPixels_ready && bufferEnable);
  assign passPixels_payload_pixel = pixelsIn_s2mPipe_m2sPipe_payload_pixel;
  assign passPixels_payload_frameStart = pixelsIn_s2mPipe_m2sPipe_payload_frameStart;
  assign passPixels_payload_rowEnd = pixelsIn_s2mPipe_m2sPipe_payload_rowEnd;
  assign passPixels_payload_inpValid = pixelsIn_s2mPipe_m2sPipe_payload_inpValid;
  assign passPixels_ready = 1'b1;
  assign passPixels_fire = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart3_l226 = ((CICC1851_when_SuperResolutionPart3_l226 == CICC1851_when_SuperResolutionPart3_l226_1) && passPixels_fire);
  assign passPixels_fire_1 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart3_l227 = (((CICC1851_when_SuperResolutionPart3_l227 == CICC1851_when_SuperResolutionPart3_l227_1) && bufferReachRowEnd) && passPixels_fire_1);
  assign passPixels_fire_2 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart3_l230 = (passPixels_payload_rowEnd && passPixels_fire_2);
  assign passPixels_fire_3 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart3_l243 = (passPixels_payload_rowEnd && passPixels_fire_3);
  assign when_SuperResolutionPart3_l244 = (bufferSwitch == 2'b10);
  assign passPixels_fire_4 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart3_l251 = (((12'h002 <= bufferRowCount_value) && passPixels_payload_rowEnd) && passPixels_fire_4);
  assign when_SuperResolutionPart3_l255 = (bufferReachFinalRow && bufferReachRowEnd);
  assign passPixels_fire_5 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart3_l262 = (passPixels_payload_frameStart && passPixels_fire_5);
  assign pixelsOut_fire = (pixelsOut_valid && pixelsOut_ready);
  assign when_SuperResolutionPart3_l270 = ((CICC1851_when_SuperResolutionPart3_l270 == CICC1851_when_SuperResolutionPart3_l270_1) && pixelsOut_fire);
  assign pixelsOut_fire_1 = (pixelsOut_valid && pixelsOut_ready);
  assign when_SuperResolutionPart3_l271 = (((CICC1851_when_SuperResolutionPart3_l271 == CICC1851_when_SuperResolutionPart3_l271_1) && alreadyReachRowEnd) && pixelsOut_fire_1);
  assign pixelsOut_fire_2 = (pixelsOut_valid && pixelsOut_ready);
  assign pixelsOut_fire_3 = (pixelsOut_valid && pixelsOut_ready);
  assign when_SuperResolutionPart3_l282 = ((alreadyReachFinalRow && alreadyReachRowEnd) && pixelsOut_fire_3);
  assign passPixels_fire_6 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_7 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_8 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_9 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_10 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_11 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_12 = (passPixels_valid && passPixels_ready);
  assign mainPixelAddrOneStream_ready = (! mainPixelAddrOneStream_rValid);
  assign mainPixelAddrOneStream_s2mPipe_valid = (mainPixelAddrOneStream_valid || mainPixelAddrOneStream_rValid);
  assign mainPixelAddrOneStream_s2mPipe_payload = (mainPixelAddrOneStream_rValid ? mainPixelAddrOneStream_rData : mainPixelAddrOneStream_payload);
  always @(*) begin
    mainPixelAddrOneStream_s2mPipe_ready = mainPixelAddrOneStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_1) begin
      mainPixelAddrOneStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_1 = (! mainPixelAddrOneStream_s2mPipe_m2sPipe_valid);
  assign mainPixelAddrOneStream_s2mPipe_m2sPipe_valid = mainPixelAddrOneStream_s2mPipe_rValid;
  assign mainPixelAddrOneStream_s2mPipe_m2sPipe_payload = mainPixelAddrOneStream_s2mPipe_rData;
  assign mainPixelAddrOneStream_s2mPipe_m2sPipe_ready = ((! CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready) || CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready = CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_mainOnePixelStream_payload = CICC1851_lineBufferOne_port1;
  assign CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_1 = readStage_mainOnePixelStream_ready;
    if(when_Stream_l368_2) begin
      CICC1851_1 = 1'b1;
    end
  end

  assign when_Stream_l368_2 = (! readStage_mainOnePixelStream_valid);
  assign readStage_mainOnePixelStream_valid = CICC1851_readStage_mainOnePixelStream_valid;
  assign readStage_mainOnePixelStream_payload = CICC1851_readStage_mainOnePixelStream_payload_2;
  assign counterPixelAddrOneStream_ready = (! counterPixelAddrOneStream_rValid);
  assign counterPixelAddrOneStream_s2mPipe_valid = (counterPixelAddrOneStream_valid || counterPixelAddrOneStream_rValid);
  assign counterPixelAddrOneStream_s2mPipe_payload = (counterPixelAddrOneStream_rValid ? counterPixelAddrOneStream_rData : counterPixelAddrOneStream_payload);
  always @(*) begin
    counterPixelAddrOneStream_s2mPipe_ready = counterPixelAddrOneStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_3) begin
      counterPixelAddrOneStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_3 = (! counterPixelAddrOneStream_s2mPipe_m2sPipe_valid);
  assign counterPixelAddrOneStream_s2mPipe_m2sPipe_valid = counterPixelAddrOneStream_s2mPipe_rValid;
  assign counterPixelAddrOneStream_s2mPipe_m2sPipe_payload = counterPixelAddrOneStream_s2mPipe_rData;
  assign counterPixelAddrOneStream_s2mPipe_m2sPipe_ready = ((! CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready) || CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready = CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_counterOnePixelStream_payload = CICC1851_lineBufferOne_port2;
  assign CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_2 = readStage_counterOnePixelStream_ready;
    if(when_Stream_l368_4) begin
      CICC1851_2 = 1'b1;
    end
  end

  assign when_Stream_l368_4 = (! readStage_counterOnePixelStream_valid);
  assign readStage_counterOnePixelStream_valid = CICC1851_readStage_counterOnePixelStream_valid;
  assign readStage_counterOnePixelStream_payload = CICC1851_readStage_counterOnePixelStream_payload_2;
  assign mainPixelAddrTwoStream_ready = (! mainPixelAddrTwoStream_rValid);
  assign mainPixelAddrTwoStream_s2mPipe_valid = (mainPixelAddrTwoStream_valid || mainPixelAddrTwoStream_rValid);
  assign mainPixelAddrTwoStream_s2mPipe_payload = (mainPixelAddrTwoStream_rValid ? mainPixelAddrTwoStream_rData : mainPixelAddrTwoStream_payload);
  always @(*) begin
    mainPixelAddrTwoStream_s2mPipe_ready = mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_5) begin
      mainPixelAddrTwoStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_5 = (! mainPixelAddrTwoStream_s2mPipe_m2sPipe_valid);
  assign mainPixelAddrTwoStream_s2mPipe_m2sPipe_valid = mainPixelAddrTwoStream_s2mPipe_rValid;
  assign mainPixelAddrTwoStream_s2mPipe_m2sPipe_payload = mainPixelAddrTwoStream_s2mPipe_rData;
  assign mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready = ((! CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready) || CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready = CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_mainTwoPixelStream_payload = CICC1851_lineBufferTwo_port1;
  assign CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_3 = readStage_mainTwoPixelStream_ready;
    if(when_Stream_l368_6) begin
      CICC1851_3 = 1'b1;
    end
  end

  assign when_Stream_l368_6 = (! readStage_mainTwoPixelStream_valid);
  assign readStage_mainTwoPixelStream_valid = CICC1851_readStage_mainTwoPixelStream_valid;
  assign readStage_mainTwoPixelStream_payload = CICC1851_readStage_mainTwoPixelStream_payload_2;
  assign counterPixelAddrTwoStream_ready = (! counterPixelAddrTwoStream_rValid);
  assign counterPixelAddrTwoStream_s2mPipe_valid = (counterPixelAddrTwoStream_valid || counterPixelAddrTwoStream_rValid);
  assign counterPixelAddrTwoStream_s2mPipe_payload = (counterPixelAddrTwoStream_rValid ? counterPixelAddrTwoStream_rData : counterPixelAddrTwoStream_payload);
  always @(*) begin
    counterPixelAddrTwoStream_s2mPipe_ready = counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_7) begin
      counterPixelAddrTwoStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_7 = (! counterPixelAddrTwoStream_s2mPipe_m2sPipe_valid);
  assign counterPixelAddrTwoStream_s2mPipe_m2sPipe_valid = counterPixelAddrTwoStream_s2mPipe_rValid;
  assign counterPixelAddrTwoStream_s2mPipe_m2sPipe_payload = counterPixelAddrTwoStream_s2mPipe_rData;
  assign counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready = ((! CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready) || CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready = CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_counterTwoPixelStream_payload = CICC1851_lineBufferTwo_port2;
  assign CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_4 = readStage_counterTwoPixelStream_ready;
    if(when_Stream_l368_8) begin
      CICC1851_4 = 1'b1;
    end
  end

  assign when_Stream_l368_8 = (! readStage_counterTwoPixelStream_valid);
  assign readStage_counterTwoPixelStream_valid = CICC1851_readStage_counterTwoPixelStream_valid;
  assign readStage_counterTwoPixelStream_payload = CICC1851_readStage_counterTwoPixelStream_payload_2;
  assign mainPixelAddrThreeStream_ready = (! mainPixelAddrThreeStream_rValid);
  assign mainPixelAddrThreeStream_s2mPipe_valid = (mainPixelAddrThreeStream_valid || mainPixelAddrThreeStream_rValid);
  assign mainPixelAddrThreeStream_s2mPipe_payload = (mainPixelAddrThreeStream_rValid ? mainPixelAddrThreeStream_rData : mainPixelAddrThreeStream_payload);
  always @(*) begin
    mainPixelAddrThreeStream_s2mPipe_ready = mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_9) begin
      mainPixelAddrThreeStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_9 = (! mainPixelAddrThreeStream_s2mPipe_m2sPipe_valid);
  assign mainPixelAddrThreeStream_s2mPipe_m2sPipe_valid = mainPixelAddrThreeStream_s2mPipe_rValid;
  assign mainPixelAddrThreeStream_s2mPipe_m2sPipe_payload = mainPixelAddrThreeStream_s2mPipe_rData;
  assign mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready = ((! CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready) || CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready = CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_mainThreePixelStream_payload = CICC1851_lineBufferThree_port1;
  assign CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_5 = readStage_mainThreePixelStream_ready;
    if(when_Stream_l368_10) begin
      CICC1851_5 = 1'b1;
    end
  end

  assign when_Stream_l368_10 = (! readStage_mainThreePixelStream_valid);
  assign readStage_mainThreePixelStream_valid = CICC1851_readStage_mainThreePixelStream_valid;
  assign readStage_mainThreePixelStream_payload = CICC1851_readStage_mainThreePixelStream_payload_2;
  assign counterPixelAddrThreeStream_ready = (! counterPixelAddrThreeStream_rValid);
  assign counterPixelAddrThreeStream_s2mPipe_valid = (counterPixelAddrThreeStream_valid || counterPixelAddrThreeStream_rValid);
  assign counterPixelAddrThreeStream_s2mPipe_payload = (counterPixelAddrThreeStream_rValid ? counterPixelAddrThreeStream_rData : counterPixelAddrThreeStream_payload);
  always @(*) begin
    counterPixelAddrThreeStream_s2mPipe_ready = counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_11) begin
      counterPixelAddrThreeStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_11 = (! counterPixelAddrThreeStream_s2mPipe_m2sPipe_valid);
  assign counterPixelAddrThreeStream_s2mPipe_m2sPipe_valid = counterPixelAddrThreeStream_s2mPipe_rValid;
  assign counterPixelAddrThreeStream_s2mPipe_m2sPipe_payload = counterPixelAddrThreeStream_s2mPipe_rData;
  assign counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready = ((! CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready) || CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready = CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_counterThreePixelStream_payload = CICC1851_lineBufferThree_port2;
  assign CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_6 = readStage_counterThreePixelStream_ready;
    if(when_Stream_l368_12) begin
      CICC1851_6 = 1'b1;
    end
  end

  assign when_Stream_l368_12 = (! readStage_counterThreePixelStream_valid);
  assign readStage_counterThreePixelStream_valid = CICC1851_readStage_counterThreePixelStream_valid;
  assign readStage_counterThreePixelStream_payload = CICC1851_readStage_counterThreePixelStream_payload_2;
  assign mainValidAddrOneStream_ready = (! mainValidAddrOneStream_rValid);
  assign mainValidAddrOneStream_s2mPipe_valid = (mainValidAddrOneStream_valid || mainValidAddrOneStream_rValid);
  assign mainValidAddrOneStream_s2mPipe_payload = (mainValidAddrOneStream_rValid ? mainValidAddrOneStream_rData : mainValidAddrOneStream_payload);
  always @(*) begin
    mainValidAddrOneStream_s2mPipe_ready = mainValidAddrOneStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_13) begin
      mainValidAddrOneStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_13 = (! mainValidAddrOneStream_s2mPipe_m2sPipe_valid);
  assign mainValidAddrOneStream_s2mPipe_m2sPipe_valid = mainValidAddrOneStream_s2mPipe_rValid;
  assign mainValidAddrOneStream_s2mPipe_m2sPipe_payload = mainValidAddrOneStream_s2mPipe_rData;
  assign mainValidAddrOneStream_s2mPipe_m2sPipe_ready = ((! CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready) || CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready = CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_mainOneValidStream_payload = CICC1851_validBufferOne_port1[0];
  assign CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_7 = readStage_mainOneValidStream_ready;
    if(when_Stream_l368_14) begin
      CICC1851_7 = 1'b1;
    end
  end

  assign when_Stream_l368_14 = (! readStage_mainOneValidStream_valid);
  assign readStage_mainOneValidStream_valid = CICC1851_readStage_mainOneValidStream_valid;
  assign readStage_mainOneValidStream_payload = CICC1851_readStage_mainOneValidStream_payload_2;
  assign counterValidAddrOneStream_ready = (! counterValidAddrOneStream_rValid);
  assign counterValidAddrOneStream_s2mPipe_valid = (counterValidAddrOneStream_valid || counterValidAddrOneStream_rValid);
  assign counterValidAddrOneStream_s2mPipe_payload = (counterValidAddrOneStream_rValid ? counterValidAddrOneStream_rData : counterValidAddrOneStream_payload);
  always @(*) begin
    counterValidAddrOneStream_s2mPipe_ready = counterValidAddrOneStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_15) begin
      counterValidAddrOneStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_15 = (! counterValidAddrOneStream_s2mPipe_m2sPipe_valid);
  assign counterValidAddrOneStream_s2mPipe_m2sPipe_valid = counterValidAddrOneStream_s2mPipe_rValid;
  assign counterValidAddrOneStream_s2mPipe_m2sPipe_payload = counterValidAddrOneStream_s2mPipe_rData;
  assign counterValidAddrOneStream_s2mPipe_m2sPipe_ready = ((! CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready) || CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready = CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_counterOneValidStream_payload = CICC1851_validBufferOne_port2[0];
  assign CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_8 = readStage_counterOneValidStream_ready;
    if(when_Stream_l368_16) begin
      CICC1851_8 = 1'b1;
    end
  end

  assign when_Stream_l368_16 = (! readStage_counterOneValidStream_valid);
  assign readStage_counterOneValidStream_valid = CICC1851_readStage_counterOneValidStream_valid;
  assign readStage_counterOneValidStream_payload = CICC1851_readStage_counterOneValidStream_payload_2;
  assign mainValidAddrTwoStream_ready = (! mainValidAddrTwoStream_rValid);
  assign mainValidAddrTwoStream_s2mPipe_valid = (mainValidAddrTwoStream_valid || mainValidAddrTwoStream_rValid);
  assign mainValidAddrTwoStream_s2mPipe_payload = (mainValidAddrTwoStream_rValid ? mainValidAddrTwoStream_rData : mainValidAddrTwoStream_payload);
  always @(*) begin
    mainValidAddrTwoStream_s2mPipe_ready = mainValidAddrTwoStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_17) begin
      mainValidAddrTwoStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_17 = (! mainValidAddrTwoStream_s2mPipe_m2sPipe_valid);
  assign mainValidAddrTwoStream_s2mPipe_m2sPipe_valid = mainValidAddrTwoStream_s2mPipe_rValid;
  assign mainValidAddrTwoStream_s2mPipe_m2sPipe_payload = mainValidAddrTwoStream_s2mPipe_rData;
  assign mainValidAddrTwoStream_s2mPipe_m2sPipe_ready = ((! CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready) || CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready = CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_mainTwoValidStream_payload = CICC1851_validBufferTwo_port1[0];
  assign CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_9 = readStage_mainTwoValidStream_ready;
    if(when_Stream_l368_18) begin
      CICC1851_9 = 1'b1;
    end
  end

  assign when_Stream_l368_18 = (! readStage_mainTwoValidStream_valid);
  assign readStage_mainTwoValidStream_valid = CICC1851_readStage_mainTwoValidStream_valid;
  assign readStage_mainTwoValidStream_payload = CICC1851_readStage_mainTwoValidStream_payload_2;
  assign counterValidAddrTwoStream_ready = (! counterValidAddrTwoStream_rValid);
  assign counterValidAddrTwoStream_s2mPipe_valid = (counterValidAddrTwoStream_valid || counterValidAddrTwoStream_rValid);
  assign counterValidAddrTwoStream_s2mPipe_payload = (counterValidAddrTwoStream_rValid ? counterValidAddrTwoStream_rData : counterValidAddrTwoStream_payload);
  always @(*) begin
    counterValidAddrTwoStream_s2mPipe_ready = counterValidAddrTwoStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_19) begin
      counterValidAddrTwoStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_19 = (! counterValidAddrTwoStream_s2mPipe_m2sPipe_valid);
  assign counterValidAddrTwoStream_s2mPipe_m2sPipe_valid = counterValidAddrTwoStream_s2mPipe_rValid;
  assign counterValidAddrTwoStream_s2mPipe_m2sPipe_payload = counterValidAddrTwoStream_s2mPipe_rData;
  assign counterValidAddrTwoStream_s2mPipe_m2sPipe_ready = ((! CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready) || CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready = CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_counterTwoValidStream_payload = CICC1851_validBufferTwo_port2[0];
  assign CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_10 = readStage_counterTwoValidStream_ready;
    if(when_Stream_l368_20) begin
      CICC1851_10 = 1'b1;
    end
  end

  assign when_Stream_l368_20 = (! readStage_counterTwoValidStream_valid);
  assign readStage_counterTwoValidStream_valid = CICC1851_readStage_counterTwoValidStream_valid;
  assign readStage_counterTwoValidStream_payload = CICC1851_readStage_counterTwoValidStream_payload_2;
  assign mainValidAddrThreeStream_ready = (! mainValidAddrThreeStream_rValid);
  assign mainValidAddrThreeStream_s2mPipe_valid = (mainValidAddrThreeStream_valid || mainValidAddrThreeStream_rValid);
  assign mainValidAddrThreeStream_s2mPipe_payload = (mainValidAddrThreeStream_rValid ? mainValidAddrThreeStream_rData : mainValidAddrThreeStream_payload);
  always @(*) begin
    mainValidAddrThreeStream_s2mPipe_ready = mainValidAddrThreeStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_21) begin
      mainValidAddrThreeStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_21 = (! mainValidAddrThreeStream_s2mPipe_m2sPipe_valid);
  assign mainValidAddrThreeStream_s2mPipe_m2sPipe_valid = mainValidAddrThreeStream_s2mPipe_rValid;
  assign mainValidAddrThreeStream_s2mPipe_m2sPipe_payload = mainValidAddrThreeStream_s2mPipe_rData;
  assign mainValidAddrThreeStream_s2mPipe_m2sPipe_ready = ((! CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready) || CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready = CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_mainThreeValidStream_payload = CICC1851_validBufferThree_port1[0];
  assign CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_11 = readStage_mainThreeValidStream_ready;
    if(when_Stream_l368_22) begin
      CICC1851_11 = 1'b1;
    end
  end

  assign when_Stream_l368_22 = (! readStage_mainThreeValidStream_valid);
  assign readStage_mainThreeValidStream_valid = CICC1851_readStage_mainThreeValidStream_valid;
  assign readStage_mainThreeValidStream_payload = CICC1851_readStage_mainThreeValidStream_payload_2;
  assign counterValidAddrThreeStream_ready = (! counterValidAddrThreeStream_rValid);
  assign counterValidAddrThreeStream_s2mPipe_valid = (counterValidAddrThreeStream_valid || counterValidAddrThreeStream_rValid);
  assign counterValidAddrThreeStream_s2mPipe_payload = (counterValidAddrThreeStream_rValid ? counterValidAddrThreeStream_rData : counterValidAddrThreeStream_payload);
  always @(*) begin
    counterValidAddrThreeStream_s2mPipe_ready = counterValidAddrThreeStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_23) begin
      counterValidAddrThreeStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_23 = (! counterValidAddrThreeStream_s2mPipe_m2sPipe_valid);
  assign counterValidAddrThreeStream_s2mPipe_m2sPipe_valid = counterValidAddrThreeStream_s2mPipe_rValid;
  assign counterValidAddrThreeStream_s2mPipe_m2sPipe_payload = counterValidAddrThreeStream_s2mPipe_rData;
  assign counterValidAddrThreeStream_s2mPipe_m2sPipe_ready = ((! CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready) || CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready = CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_counterThreeValidStream_payload = CICC1851_validBufferThree_port2[0];
  assign CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_12 = readStage_counterThreeValidStream_ready;
    if(when_Stream_l368_24) begin
      CICC1851_12 = 1'b1;
    end
  end

  assign when_Stream_l368_24 = (! readStage_counterThreeValidStream_valid);
  assign readStage_counterThreeValidStream_valid = CICC1851_readStage_counterThreeValidStream_valid;
  assign readStage_counterThreeValidStream_payload = CICC1851_readStage_counterThreeValidStream_payload_2;
  assign controlStream_ready = (! controlStream_rValid);
  assign controlStream_s2mPipe_valid = (controlStream_valid || controlStream_rValid);
  assign controlStream_s2mPipe_payload_frameStart = (controlStream_rValid ? controlStream_rData_frameStart : controlStream_payload_frameStart);
  assign controlStream_s2mPipe_payload_rowEnd = (controlStream_rValid ? controlStream_rData_rowEnd : controlStream_payload_rowEnd);
  assign controlStream_s2mPipe_payload_pipeValid = (controlStream_rValid ? controlStream_rData_pipeValid : controlStream_payload_pipeValid);
  assign controlStream_s2mPipe_payload_firstRow = (controlStream_rValid ? controlStream_rData_firstRow : controlStream_payload_firstRow);
  assign controlStream_s2mPipe_payload_lastRow = (controlStream_rValid ? controlStream_rData_lastRow : controlStream_payload_lastRow);
  assign controlStream_s2mPipe_payload_finalResult = (controlStream_rValid ? controlStream_rData_finalResult : controlStream_payload_finalResult);
  assign controlStream_s2mPipe_payload_mainCompare = (controlStream_rValid ? controlStream_rData_mainCompare : controlStream_payload_mainCompare);
  assign controlStream_s2mPipe_payload_counterCompare = (controlStream_rValid ? controlStream_rData_counterCompare : controlStream_payload_counterCompare);
  assign controlStream_s2mPipe_payload_horizontalCompare = (controlStream_rValid ? controlStream_rData_horizontalCompare : controlStream_payload_horizontalCompare);
  assign controlStream_s2mPipe_payload_verticalCompare = (controlStream_rValid ? controlStream_rData_verticalCompare : controlStream_payload_verticalCompare);
  assign controlStream_s2mPipe_payload_mainDiff = (controlStream_rValid ? controlStream_rData_mainDiff : controlStream_payload_mainDiff);
  assign controlStream_s2mPipe_payload_counterDiff = (controlStream_rValid ? controlStream_rData_counterDiff : controlStream_payload_counterDiff);
  assign controlStream_s2mPipe_payload_horizontalDiff = (controlStream_rValid ? controlStream_rData_horizontalDiff : controlStream_payload_horizontalDiff);
  assign controlStream_s2mPipe_payload_verticalDiff = (controlStream_rValid ? controlStream_rData_verticalDiff : controlStream_payload_verticalDiff);
  assign controlStream_s2mPipe_payload_isHorizontalMin = (controlStream_rValid ? controlStream_rData_isHorizontalMin : controlStream_payload_isHorizontalMin);
  assign controlStream_s2mPipe_payload_minDiff = (controlStream_rValid ? controlStream_rData_minDiff : controlStream_payload_minDiff);
  assign controlStream_s2mPipe_payload_currentPosition = (controlStream_rValid ? controlStream_rData_currentPosition : controlStream_payload_currentPosition);
  assign controlStream_s2mPipe_payload_nextPosition = (controlStream_rValid ? controlStream_rData_nextPosition : controlStream_payload_nextPosition);
  assign controlStream_s2mPipe_payload_horizontalDirectionValid = (controlStream_rValid ? controlStream_rData_horizontalDirectionValid : controlStream_payload_horizontalDirectionValid);
  assign controlStream_s2mPipe_payload_verticalDirectionValid = (controlStream_rValid ? controlStream_rData_verticalDirectionValid : controlStream_payload_verticalDirectionValid);
  assign controlStream_s2mPipe_payload_mainDirectionValid = (controlStream_rValid ? controlStream_rData_mainDirectionValid : controlStream_payload_mainDirectionValid);
  assign controlStream_s2mPipe_payload_counterDirectionValid = (controlStream_rValid ? controlStream_rData_counterDirectionValid : controlStream_payload_counterDirectionValid);
  assign controlStream_s2mPipe_payload_inValidMinDiff = (controlStream_rValid ? controlStream_rData_inValidMinDiff : controlStream_payload_inValidMinDiff);
  always @(*) begin
    controlStream_s2mPipe_ready = controlStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_25) begin
      controlStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_25 = (! controlStream_s2mPipe_m2sPipe_valid);
  assign controlStream_s2mPipe_m2sPipe_valid = controlStream_s2mPipe_rValid;
  assign controlStream_s2mPipe_m2sPipe_payload_frameStart = controlStream_s2mPipe_rData_frameStart;
  assign controlStream_s2mPipe_m2sPipe_payload_rowEnd = controlStream_s2mPipe_rData_rowEnd;
  assign controlStream_s2mPipe_m2sPipe_payload_pipeValid = controlStream_s2mPipe_rData_pipeValid;
  assign controlStream_s2mPipe_m2sPipe_payload_firstRow = controlStream_s2mPipe_rData_firstRow;
  assign controlStream_s2mPipe_m2sPipe_payload_lastRow = controlStream_s2mPipe_rData_lastRow;
  assign controlStream_s2mPipe_m2sPipe_payload_finalResult = controlStream_s2mPipe_rData_finalResult;
  assign controlStream_s2mPipe_m2sPipe_payload_mainCompare = controlStream_s2mPipe_rData_mainCompare;
  assign controlStream_s2mPipe_m2sPipe_payload_counterCompare = controlStream_s2mPipe_rData_counterCompare;
  assign controlStream_s2mPipe_m2sPipe_payload_horizontalCompare = controlStream_s2mPipe_rData_horizontalCompare;
  assign controlStream_s2mPipe_m2sPipe_payload_verticalCompare = controlStream_s2mPipe_rData_verticalCompare;
  assign controlStream_s2mPipe_m2sPipe_payload_mainDiff = controlStream_s2mPipe_rData_mainDiff;
  assign controlStream_s2mPipe_m2sPipe_payload_counterDiff = controlStream_s2mPipe_rData_counterDiff;
  assign controlStream_s2mPipe_m2sPipe_payload_horizontalDiff = controlStream_s2mPipe_rData_horizontalDiff;
  assign controlStream_s2mPipe_m2sPipe_payload_verticalDiff = controlStream_s2mPipe_rData_verticalDiff;
  assign controlStream_s2mPipe_m2sPipe_payload_isHorizontalMin = controlStream_s2mPipe_rData_isHorizontalMin;
  assign controlStream_s2mPipe_m2sPipe_payload_minDiff = controlStream_s2mPipe_rData_minDiff;
  assign controlStream_s2mPipe_m2sPipe_payload_currentPosition = controlStream_s2mPipe_rData_currentPosition;
  assign controlStream_s2mPipe_m2sPipe_payload_nextPosition = controlStream_s2mPipe_rData_nextPosition;
  assign controlStream_s2mPipe_m2sPipe_payload_horizontalDirectionValid = controlStream_s2mPipe_rData_horizontalDirectionValid;
  assign controlStream_s2mPipe_m2sPipe_payload_verticalDirectionValid = controlStream_s2mPipe_rData_verticalDirectionValid;
  assign controlStream_s2mPipe_m2sPipe_payload_mainDirectionValid = controlStream_s2mPipe_rData_mainDirectionValid;
  assign controlStream_s2mPipe_m2sPipe_payload_counterDirectionValid = controlStream_s2mPipe_rData_counterDirectionValid;
  assign controlStream_s2mPipe_m2sPipe_payload_inValidMinDiff = controlStream_s2mPipe_rData_inValidMinDiff;
  always @(*) begin
    controlStream_s2mPipe_m2sPipe_ready = controlStream_s2mPipe_m2sPipe_m2sPipe_ready;
    if(when_Stream_l368_26) begin
      controlStream_s2mPipe_m2sPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_26 = (! controlStream_s2mPipe_m2sPipe_m2sPipe_valid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_valid = controlStream_s2mPipe_m2sPipe_rValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_frameStart = controlStream_s2mPipe_m2sPipe_rData_frameStart;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_rowEnd = controlStream_s2mPipe_m2sPipe_rData_rowEnd;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_pipeValid = controlStream_s2mPipe_m2sPipe_rData_pipeValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_firstRow = controlStream_s2mPipe_m2sPipe_rData_firstRow;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_lastRow = controlStream_s2mPipe_m2sPipe_rData_lastRow;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_finalResult = controlStream_s2mPipe_m2sPipe_rData_finalResult;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainCompare = controlStream_s2mPipe_m2sPipe_rData_mainCompare;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterCompare = controlStream_s2mPipe_m2sPipe_rData_counterCompare;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_horizontalCompare = controlStream_s2mPipe_m2sPipe_rData_horizontalCompare;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_verticalCompare = controlStream_s2mPipe_m2sPipe_rData_verticalCompare;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDiff = controlStream_s2mPipe_m2sPipe_rData_mainDiff;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDiff = controlStream_s2mPipe_m2sPipe_rData_counterDiff;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_horizontalDiff = controlStream_s2mPipe_m2sPipe_rData_horizontalDiff;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_verticalDiff = controlStream_s2mPipe_m2sPipe_rData_verticalDiff;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_isHorizontalMin = controlStream_s2mPipe_m2sPipe_rData_isHorizontalMin;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_minDiff = controlStream_s2mPipe_m2sPipe_rData_minDiff;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_currentPosition = controlStream_s2mPipe_m2sPipe_rData_currentPosition;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_nextPosition = controlStream_s2mPipe_m2sPipe_rData_nextPosition;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_horizontalDirectionValid = controlStream_s2mPipe_m2sPipe_rData_horizontalDirectionValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_verticalDirectionValid = controlStream_s2mPipe_m2sPipe_rData_verticalDirectionValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDirectionValid = controlStream_s2mPipe_m2sPipe_rData_mainDirectionValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDirectionValid = controlStream_s2mPipe_m2sPipe_rData_counterDirectionValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_inValidMinDiff = controlStream_s2mPipe_m2sPipe_rData_inValidMinDiff;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_ready = (! controlStream_s2mPipe_m2sPipe_m2sPipe_rValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_valid = (controlStream_s2mPipe_m2sPipe_m2sPipe_valid || controlStream_s2mPipe_m2sPipe_m2sPipe_rValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_frameStart = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_frameStart : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_frameStart);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_rowEnd = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_rowEnd : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_rowEnd);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_pipeValid = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_pipeValid : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_pipeValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_firstRow = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_firstRow : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_firstRow);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_lastRow = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_lastRow : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_lastRow);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_finalResult = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_finalResult : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_finalResult);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainCompare = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainCompare : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainCompare);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterCompare = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterCompare : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterCompare);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_horizontalCompare = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_horizontalCompare : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_horizontalCompare);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_verticalCompare = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_verticalCompare : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_verticalCompare);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainDiff = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainDiff : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDiff);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterDiff = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterDiff : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDiff);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_horizontalDiff = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_horizontalDiff : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_horizontalDiff);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_verticalDiff = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_verticalDiff : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_verticalDiff);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_isHorizontalMin = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_isHorizontalMin : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_isHorizontalMin);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_minDiff = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_minDiff : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_minDiff);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_currentPosition = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_currentPosition : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_currentPosition);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_nextPosition = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_nextPosition : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_nextPosition);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_horizontalDirectionValid = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_horizontalDirectionValid : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_horizontalDirectionValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_verticalDirectionValid = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_verticalDirectionValid : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_verticalDirectionValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainDirectionValid = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainDirectionValid : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDirectionValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterDirectionValid = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterDirectionValid : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDirectionValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_inValidMinDiff = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_inValidMinDiff : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_inValidMinDiff);
  always @(*) begin
    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready = readStage_controlPipe_ready;
    if(when_Stream_l368_27) begin
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_27 = (! readStage_controlPipe_valid);
  assign readStage_controlPipe_valid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rValid;
  assign readStage_controlPipe_payload_frameStart = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_frameStart;
  assign readStage_controlPipe_payload_rowEnd = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_rowEnd;
  assign readStage_controlPipe_payload_pipeValid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_pipeValid;
  assign readStage_controlPipe_payload_firstRow = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_firstRow;
  assign readStage_controlPipe_payload_lastRow = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_lastRow;
  assign readStage_controlPipe_payload_finalResult = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_finalResult;
  assign readStage_controlPipe_payload_mainCompare = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainCompare;
  assign readStage_controlPipe_payload_counterCompare = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterCompare;
  assign readStage_controlPipe_payload_horizontalCompare = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_horizontalCompare;
  assign readStage_controlPipe_payload_verticalCompare = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_verticalCompare;
  assign readStage_controlPipe_payload_mainDiff = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainDiff;
  assign readStage_controlPipe_payload_counterDiff = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterDiff;
  assign readStage_controlPipe_payload_horizontalDiff = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_horizontalDiff;
  assign readStage_controlPipe_payload_verticalDiff = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_verticalDiff;
  assign readStage_controlPipe_payload_isHorizontalMin = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_isHorizontalMin;
  assign readStage_controlPipe_payload_minDiff = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_minDiff;
  assign readStage_controlPipe_payload_currentPosition = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_currentPosition;
  assign readStage_controlPipe_payload_nextPosition = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_nextPosition;
  assign readStage_controlPipe_payload_horizontalDirectionValid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_horizontalDirectionValid;
  assign readStage_controlPipe_payload_verticalDirectionValid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_verticalDirectionValid;
  assign readStage_controlPipe_payload_mainDirectionValid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainDirectionValid;
  assign readStage_controlPipe_payload_counterDirectionValid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterDirectionValid;
  assign readStage_controlPipe_payload_inValidMinDiff = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_inValidMinDiff;
  assign readStage_mainOnePixelStream_ready = (! readStage_mainOnePixelStream_rValid);
  assign readStage_mainOnePixelStream_s2mPipe_valid = (readStage_mainOnePixelStream_valid || readStage_mainOnePixelStream_rValid);
  assign readStage_mainOnePixelStream_s2mPipe_payload = (readStage_mainOnePixelStream_rValid ? readStage_mainOnePixelStream_rData : readStage_mainOnePixelStream_payload);
  always @(*) begin
    readStage_mainOnePixelStream_s2mPipe_ready = compareStage_mainOnePixelStream_ready;
    if(when_Stream_l368_28) begin
      readStage_mainOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_28 = (! compareStage_mainOnePixelStream_valid);
  assign compareStage_mainOnePixelStream_valid = readStage_mainOnePixelStream_s2mPipe_rValid;
  assign compareStage_mainOnePixelStream_payload = readStage_mainOnePixelStream_s2mPipe_rData;
  assign readStage_counterOnePixelStream_ready = (! readStage_counterOnePixelStream_rValid);
  assign readStage_counterOnePixelStream_s2mPipe_valid = (readStage_counterOnePixelStream_valid || readStage_counterOnePixelStream_rValid);
  assign readStage_counterOnePixelStream_s2mPipe_payload = (readStage_counterOnePixelStream_rValid ? readStage_counterOnePixelStream_rData : readStage_counterOnePixelStream_payload);
  always @(*) begin
    readStage_counterOnePixelStream_s2mPipe_ready = compareStage_counterOnePixelStream_ready;
    if(when_Stream_l368_29) begin
      readStage_counterOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_29 = (! compareStage_counterOnePixelStream_valid);
  assign compareStage_counterOnePixelStream_valid = readStage_counterOnePixelStream_s2mPipe_rValid;
  assign compareStage_counterOnePixelStream_payload = readStage_counterOnePixelStream_s2mPipe_rData;
  assign readStage_mainTwoPixelStream_ready = (! readStage_mainTwoPixelStream_rValid);
  assign readStage_mainTwoPixelStream_s2mPipe_valid = (readStage_mainTwoPixelStream_valid || readStage_mainTwoPixelStream_rValid);
  assign readStage_mainTwoPixelStream_s2mPipe_payload = (readStage_mainTwoPixelStream_rValid ? readStage_mainTwoPixelStream_rData : readStage_mainTwoPixelStream_payload);
  always @(*) begin
    readStage_mainTwoPixelStream_s2mPipe_ready = compareStage_mainTwoPixelStream_ready;
    if(when_Stream_l368_30) begin
      readStage_mainTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_30 = (! compareStage_mainTwoPixelStream_valid);
  assign compareStage_mainTwoPixelStream_valid = readStage_mainTwoPixelStream_s2mPipe_rValid;
  assign compareStage_mainTwoPixelStream_payload = readStage_mainTwoPixelStream_s2mPipe_rData;
  assign readStage_counterTwoPixelStream_ready = (! readStage_counterTwoPixelStream_rValid);
  assign readStage_counterTwoPixelStream_s2mPipe_valid = (readStage_counterTwoPixelStream_valid || readStage_counterTwoPixelStream_rValid);
  assign readStage_counterTwoPixelStream_s2mPipe_payload = (readStage_counterTwoPixelStream_rValid ? readStage_counterTwoPixelStream_rData : readStage_counterTwoPixelStream_payload);
  always @(*) begin
    readStage_counterTwoPixelStream_s2mPipe_ready = compareStage_counterTwoPixelStream_ready;
    if(when_Stream_l368_31) begin
      readStage_counterTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_31 = (! compareStage_counterTwoPixelStream_valid);
  assign compareStage_counterTwoPixelStream_valid = readStage_counterTwoPixelStream_s2mPipe_rValid;
  assign compareStage_counterTwoPixelStream_payload = readStage_counterTwoPixelStream_s2mPipe_rData;
  assign readStage_mainThreePixelStream_ready = (! readStage_mainThreePixelStream_rValid);
  assign readStage_mainThreePixelStream_s2mPipe_valid = (readStage_mainThreePixelStream_valid || readStage_mainThreePixelStream_rValid);
  assign readStage_mainThreePixelStream_s2mPipe_payload = (readStage_mainThreePixelStream_rValid ? readStage_mainThreePixelStream_rData : readStage_mainThreePixelStream_payload);
  always @(*) begin
    readStage_mainThreePixelStream_s2mPipe_ready = compareStage_mainThreePixelStream_ready;
    if(when_Stream_l368_32) begin
      readStage_mainThreePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_32 = (! compareStage_mainThreePixelStream_valid);
  assign compareStage_mainThreePixelStream_valid = readStage_mainThreePixelStream_s2mPipe_rValid;
  assign compareStage_mainThreePixelStream_payload = readStage_mainThreePixelStream_s2mPipe_rData;
  assign readStage_counterThreePixelStream_ready = (! readStage_counterThreePixelStream_rValid);
  assign readStage_counterThreePixelStream_s2mPipe_valid = (readStage_counterThreePixelStream_valid || readStage_counterThreePixelStream_rValid);
  assign readStage_counterThreePixelStream_s2mPipe_payload = (readStage_counterThreePixelStream_rValid ? readStage_counterThreePixelStream_rData : readStage_counterThreePixelStream_payload);
  always @(*) begin
    readStage_counterThreePixelStream_s2mPipe_ready = compareStage_counterThreePixelStream_ready;
    if(when_Stream_l368_33) begin
      readStage_counterThreePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_33 = (! compareStage_counterThreePixelStream_valid);
  assign compareStage_counterThreePixelStream_valid = readStage_counterThreePixelStream_s2mPipe_rValid;
  assign compareStage_counterThreePixelStream_payload = readStage_counterThreePixelStream_s2mPipe_rData;
  assign readStage_mainOneValidStream_ready = (! readStage_mainOneValidStream_rValid);
  assign readStage_mainOneValidStream_s2mPipe_valid = (readStage_mainOneValidStream_valid || readStage_mainOneValidStream_rValid);
  assign readStage_mainOneValidStream_s2mPipe_payload = (readStage_mainOneValidStream_rValid ? readStage_mainOneValidStream_rData : readStage_mainOneValidStream_payload);
  always @(*) begin
    readStage_mainOneValidStream_s2mPipe_ready = compareStage_mainOneValidStream_ready;
    if(when_Stream_l368_34) begin
      readStage_mainOneValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_34 = (! compareStage_mainOneValidStream_valid);
  assign compareStage_mainOneValidStream_valid = readStage_mainOneValidStream_s2mPipe_rValid;
  assign compareStage_mainOneValidStream_payload = readStage_mainOneValidStream_s2mPipe_rData;
  assign readStage_counterOneValidStream_ready = (! readStage_counterOneValidStream_rValid);
  assign readStage_counterOneValidStream_s2mPipe_valid = (readStage_counterOneValidStream_valid || readStage_counterOneValidStream_rValid);
  assign readStage_counterOneValidStream_s2mPipe_payload = (readStage_counterOneValidStream_rValid ? readStage_counterOneValidStream_rData : readStage_counterOneValidStream_payload);
  always @(*) begin
    readStage_counterOneValidStream_s2mPipe_ready = compareStage_counterOneValidStream_ready;
    if(when_Stream_l368_35) begin
      readStage_counterOneValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_35 = (! compareStage_counterOneValidStream_valid);
  assign compareStage_counterOneValidStream_valid = readStage_counterOneValidStream_s2mPipe_rValid;
  assign compareStage_counterOneValidStream_payload = readStage_counterOneValidStream_s2mPipe_rData;
  assign readStage_mainTwoValidStream_ready = (! readStage_mainTwoValidStream_rValid);
  assign readStage_mainTwoValidStream_s2mPipe_valid = (readStage_mainTwoValidStream_valid || readStage_mainTwoValidStream_rValid);
  assign readStage_mainTwoValidStream_s2mPipe_payload = (readStage_mainTwoValidStream_rValid ? readStage_mainTwoValidStream_rData : readStage_mainTwoValidStream_payload);
  always @(*) begin
    readStage_mainTwoValidStream_s2mPipe_ready = compareStage_mainTwoValidStream_ready;
    if(when_Stream_l368_36) begin
      readStage_mainTwoValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_36 = (! compareStage_mainTwoValidStream_valid);
  assign compareStage_mainTwoValidStream_valid = readStage_mainTwoValidStream_s2mPipe_rValid;
  assign compareStage_mainTwoValidStream_payload = readStage_mainTwoValidStream_s2mPipe_rData;
  assign readStage_counterTwoValidStream_ready = (! readStage_counterTwoValidStream_rValid);
  assign readStage_counterTwoValidStream_s2mPipe_valid = (readStage_counterTwoValidStream_valid || readStage_counterTwoValidStream_rValid);
  assign readStage_counterTwoValidStream_s2mPipe_payload = (readStage_counterTwoValidStream_rValid ? readStage_counterTwoValidStream_rData : readStage_counterTwoValidStream_payload);
  always @(*) begin
    readStage_counterTwoValidStream_s2mPipe_ready = compareStage_counterTwoValidStream_ready;
    if(when_Stream_l368_37) begin
      readStage_counterTwoValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_37 = (! compareStage_counterTwoValidStream_valid);
  assign compareStage_counterTwoValidStream_valid = readStage_counterTwoValidStream_s2mPipe_rValid;
  assign compareStage_counterTwoValidStream_payload = readStage_counterTwoValidStream_s2mPipe_rData;
  assign readStage_mainThreeValidStream_ready = (! readStage_mainThreeValidStream_rValid);
  assign readStage_mainThreeValidStream_s2mPipe_valid = (readStage_mainThreeValidStream_valid || readStage_mainThreeValidStream_rValid);
  assign readStage_mainThreeValidStream_s2mPipe_payload = (readStage_mainThreeValidStream_rValid ? readStage_mainThreeValidStream_rData : readStage_mainThreeValidStream_payload);
  always @(*) begin
    readStage_mainThreeValidStream_s2mPipe_ready = compareStage_mainThreeValidStream_ready;
    if(when_Stream_l368_38) begin
      readStage_mainThreeValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_38 = (! compareStage_mainThreeValidStream_valid);
  assign compareStage_mainThreeValidStream_valid = readStage_mainThreeValidStream_s2mPipe_rValid;
  assign compareStage_mainThreeValidStream_payload = readStage_mainThreeValidStream_s2mPipe_rData;
  assign readStage_counterThreeValidStream_ready = (! readStage_counterThreeValidStream_rValid);
  assign readStage_counterThreeValidStream_s2mPipe_valid = (readStage_counterThreeValidStream_valid || readStage_counterThreeValidStream_rValid);
  assign readStage_counterThreeValidStream_s2mPipe_payload = (readStage_counterThreeValidStream_rValid ? readStage_counterThreeValidStream_rData : readStage_counterThreeValidStream_payload);
  always @(*) begin
    readStage_counterThreeValidStream_s2mPipe_ready = compareStage_counterThreeValidStream_ready;
    if(when_Stream_l368_39) begin
      readStage_counterThreeValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_39 = (! compareStage_counterThreeValidStream_valid);
  assign compareStage_counterThreeValidStream_valid = readStage_counterThreeValidStream_s2mPipe_rValid;
  assign compareStage_counterThreeValidStream_payload = readStage_counterThreeValidStream_s2mPipe_rData;
  always @(*) begin
    CICC1851_readStage_controlPipe_translated_payload_mainCompare = readStage_controlPipe_payload_mainCompare;
    if(!readStage_controlPipe_payload_finalResult) begin
      if(when_SuperResolutionPart3_l415) begin
        if(when_SuperResolutionPart3_l422) begin
          if(readStage_controlPipe_payload_firstRow) begin
            if(when_SuperResolutionPart3_l432) begin
              CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l449) begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l463) begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
              end
            end
          end
        end else begin
          if(readStage_controlPipe_payload_lastRow) begin
            if(when_SuperResolutionPart3_l477) begin
              CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
            end
          end else begin
            if(when_SuperResolutionPart3_l490) begin
              CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
            end
          end
        end
      end else begin
        if(when_SuperResolutionPart3_l496) begin
          if(when_SuperResolutionPart3_l502) begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l511) begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l524) begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
              end
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l539) begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l552) begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
              end
            end
          end
        end else begin
          if(when_SuperResolutionPart3_l564) begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l573) begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l586) begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
              end
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l601) begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l614) begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
              end
            end
          end
        end
      end
    end
  end

  always @(*) begin
    CICC1851_readStage_controlPipe_translated_payload_counterCompare = readStage_controlPipe_payload_counterCompare;
    if(!readStage_controlPipe_payload_finalResult) begin
      if(when_SuperResolutionPart3_l415) begin
        if(when_SuperResolutionPart3_l422) begin
          if(readStage_controlPipe_payload_firstRow) begin
            if(when_SuperResolutionPart3_l432) begin
              CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l449) begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l465) begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
              end
            end
          end
        end else begin
          if(readStage_controlPipe_payload_lastRow) begin
            if(when_SuperResolutionPart3_l477) begin
              CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
            end
          end else begin
            if(when_SuperResolutionPart3_l492) begin
              CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
            end
          end
        end
      end else begin
        if(when_SuperResolutionPart3_l496) begin
          if(when_SuperResolutionPart3_l502) begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l511) begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l526) begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
              end
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l539) begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l554) begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
              end
            end
          end
        end else begin
          if(when_SuperResolutionPart3_l564) begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l573) begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l588) begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
              end
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l601) begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l616) begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
              end
            end
          end
        end
      end
    end
  end

  always @(*) begin
    CICC1851_readStage_controlPipe_translated_payload_horizontalCompare = readStage_controlPipe_payload_horizontalCompare;
    if(!readStage_controlPipe_payload_finalResult) begin
      if(when_SuperResolutionPart3_l415) begin
        if(when_SuperResolutionPart3_l419) begin
          CICC1851_readStage_controlPipe_translated_payload_horizontalCompare = 1'b1;
        end else begin
          CICC1851_readStage_controlPipe_translated_payload_horizontalCompare = 1'b0;
        end
      end else begin
        if(when_SuperResolutionPart3_l496) begin
          if(when_SuperResolutionPart3_l500) begin
            CICC1851_readStage_controlPipe_translated_payload_horizontalCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_horizontalCompare = 1'b0;
          end
        end else begin
          if(when_SuperResolutionPart3_l562) begin
            CICC1851_readStage_controlPipe_translated_payload_horizontalCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_horizontalCompare = 1'b0;
          end
        end
      end
    end
  end

  always @(*) begin
    CICC1851_readStage_controlPipe_translated_payload_verticalCompare = readStage_controlPipe_payload_verticalCompare;
    if(readStage_controlPipe_payload_finalResult) begin
      if(when_SuperResolutionPart3_l342) begin
        CICC1851_readStage_controlPipe_translated_payload_verticalCompare = 1'b1;
      end else begin
        if(when_SuperResolutionPart3_l344) begin
          if(when_SuperResolutionPart3_l345) begin
            CICC1851_readStage_controlPipe_translated_payload_verticalCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_verticalCompare = 1'b0;
          end
        end else begin
          if(when_SuperResolutionPart3_l347) begin
            if(when_SuperResolutionPart3_l348) begin
              CICC1851_readStage_controlPipe_translated_payload_verticalCompare = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_verticalCompare = 1'b0;
            end
          end else begin
            if(when_SuperResolutionPart3_l351) begin
              CICC1851_readStage_controlPipe_translated_payload_verticalCompare = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_verticalCompare = 1'b0;
            end
          end
        end
      end
    end
  end

  always @(*) begin
    CICC1851_readStage_controlPipe_translated_payload_horizontalDirectionValid = readStage_controlPipe_payload_horizontalDirectionValid;
    if(!readStage_controlPipe_payload_finalResult) begin
      if(when_SuperResolutionPart3_l415) begin
        if(when_SuperResolutionPart3_l416) begin
          CICC1851_readStage_controlPipe_translated_payload_horizontalDirectionValid = 1'b1;
        end else begin
          CICC1851_readStage_controlPipe_translated_payload_horizontalDirectionValid = 1'b0;
        end
      end else begin
        if(when_SuperResolutionPart3_l496) begin
          if(when_SuperResolutionPart3_l497) begin
            CICC1851_readStage_controlPipe_translated_payload_horizontalDirectionValid = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_horizontalDirectionValid = 1'b0;
          end
        end else begin
          if(when_SuperResolutionPart3_l559) begin
            CICC1851_readStage_controlPipe_translated_payload_horizontalDirectionValid = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_horizontalDirectionValid = 1'b0;
          end
        end
      end
    end
  end

  always @(*) begin
    CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = readStage_controlPipe_payload_verticalDirectionValid;
    if(readStage_controlPipe_payload_finalResult) begin
      if(when_SuperResolutionPart3_l356) begin
        if(when_SuperResolutionPart3_l357) begin
          if(readStage_controlPipe_payload_firstRow) begin
            if(readStage_mainTwoValidStream_payload) begin
              CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b0;
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(readStage_mainThreeValidStream_payload) begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l365) begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b0;
              end
            end
          end
        end else begin
          if(readStage_controlPipe_payload_lastRow) begin
            if(readStage_mainTwoValidStream_payload) begin
              CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b0;
            end
          end else begin
            if(when_SuperResolutionPart3_l373) begin
              CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b0;
            end
          end
        end
      end else begin
        if(when_SuperResolutionPart3_l377) begin
          if(when_SuperResolutionPart3_l378) begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(readStage_mainThreeValidStream_payload) begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l383) begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b0;
              end
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(readStage_mainOneValidStream_payload) begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l391) begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b0;
              end
            end
          end
        end else begin
          if(when_SuperResolutionPart3_l396) begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(readStage_mainTwoValidStream_payload) begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l401) begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b0;
              end
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(readStage_mainOneValidStream_payload) begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l409) begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b0;
              end
            end
          end
        end
      end
    end
  end

  always @(*) begin
    CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = readStage_controlPipe_payload_mainDirectionValid;
    if(!readStage_controlPipe_payload_finalResult) begin
      if(when_SuperResolutionPart3_l415) begin
        if(when_SuperResolutionPart3_l422) begin
          if(readStage_controlPipe_payload_firstRow) begin
            if(when_SuperResolutionPart3_l424) begin
              CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b0;
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l441) begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l458) begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b0;
              end
            end
          end
        end else begin
          if(readStage_controlPipe_payload_lastRow) begin
            if(when_SuperResolutionPart3_l470) begin
              CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b0;
            end
          end else begin
            if(when_SuperResolutionPart3_l485) begin
              CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b0;
            end
          end
        end
      end else begin
        if(when_SuperResolutionPart3_l496) begin
          if(when_SuperResolutionPart3_l502) begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l504) begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l519) begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b0;
              end
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l531) begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l547) begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b0;
              end
            end
          end
        end else begin
          if(when_SuperResolutionPart3_l564) begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l566) begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l581) begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b0;
              end
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l593) begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l609) begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b0;
              end
            end
          end
        end
      end
    end
  end

  always @(*) begin
    CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = readStage_controlPipe_payload_counterDirectionValid;
    if(!readStage_controlPipe_payload_finalResult) begin
      if(when_SuperResolutionPart3_l415) begin
        if(when_SuperResolutionPart3_l422) begin
          if(readStage_controlPipe_payload_firstRow) begin
            if(when_SuperResolutionPart3_l424) begin
              CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b0;
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l441) begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l460) begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b0;
              end
            end
          end
        end else begin
          if(readStage_controlPipe_payload_lastRow) begin
            if(when_SuperResolutionPart3_l470) begin
              CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b0;
            end
          end else begin
            if(when_SuperResolutionPart3_l487) begin
              CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b0;
            end
          end
        end
      end else begin
        if(when_SuperResolutionPart3_l496) begin
          if(when_SuperResolutionPart3_l502) begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l504) begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l521) begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b0;
              end
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l531) begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l549) begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b0;
              end
            end
          end
        end else begin
          if(when_SuperResolutionPart3_l564) begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l566) begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l583) begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b0;
              end
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l593) begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l611) begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b0;
              end
            end
          end
        end
      end
    end
  end

  assign when_SuperResolutionPart3_l342 = (readStage_controlPipe_payload_firstRow || readStage_controlPipe_payload_lastRow);
  assign when_SuperResolutionPart3_l344 = (readStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l345 = (readStage_mainThreePixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart3_l348 = (readStage_mainThreePixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart3_l351 = (readStage_mainTwoPixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart3_l347 = (readStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l356 = (readStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l357 = (readStage_controlPipe_payload_nextPosition == 2'b01);
  assign when_SuperResolutionPart3_l365 = (readStage_mainTwoValidStream_payload && readStage_mainThreeValidStream_payload);
  assign when_SuperResolutionPart3_l373 = (readStage_mainTwoValidStream_payload && readStage_mainThreeValidStream_payload);
  assign when_SuperResolutionPart3_l378 = (readStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l383 = (readStage_mainOneValidStream_payload && readStage_mainThreeValidStream_payload);
  assign when_SuperResolutionPart3_l391 = (readStage_mainOneValidStream_payload && readStage_mainThreeValidStream_payload);
  assign when_SuperResolutionPart3_l396 = (readStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l401 = (readStage_mainOneValidStream_payload && readStage_mainTwoValidStream_payload);
  assign when_SuperResolutionPart3_l409 = (readStage_mainOneValidStream_payload && readStage_mainTwoValidStream_payload);
  assign when_SuperResolutionPart3_l377 = (readStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l415 = (readStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l416 = (readStage_mainOneValidStream_payload && readStage_counterOneValidStream_payload);
  assign when_SuperResolutionPart3_l419 = (readStage_counterOnePixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart3_l422 = (readStage_controlPipe_payload_nextPosition == 2'b01);
  assign when_SuperResolutionPart3_l424 = (readStage_mainTwoValidStream_payload && readStage_counterTwoValidStream_payload);
  assign when_SuperResolutionPart3_l432 = (readStage_counterTwoPixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart3_l441 = (readStage_mainThreeValidStream_payload && readStage_counterThreeValidStream_payload);
  assign when_SuperResolutionPart3_l449 = (readStage_counterThreePixelStream_payload <= readStage_mainThreePixelStream_payload);
  assign when_SuperResolutionPart3_l458 = (readStage_mainThreeValidStream_payload && readStage_counterTwoValidStream_payload);
  assign when_SuperResolutionPart3_l460 = (readStage_mainTwoValidStream_payload && readStage_counterThreeValidStream_payload);
  assign when_SuperResolutionPart3_l463 = (readStage_counterTwoPixelStream_payload <= readStage_mainThreePixelStream_payload);
  assign when_SuperResolutionPart3_l465 = (readStage_counterThreePixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart3_l470 = (readStage_mainTwoValidStream_payload && readStage_counterTwoValidStream_payload);
  assign when_SuperResolutionPart3_l477 = (readStage_counterTwoPixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart3_l485 = (readStage_mainTwoValidStream_payload && readStage_counterThreeValidStream_payload);
  assign when_SuperResolutionPart3_l487 = (readStage_mainThreeValidStream_payload && readStage_counterTwoValidStream_payload);
  assign when_SuperResolutionPart3_l490 = (readStage_counterThreePixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart3_l492 = (readStage_counterTwoPixelStream_payload <= readStage_mainThreePixelStream_payload);
  assign when_SuperResolutionPart3_l497 = (readStage_mainTwoValidStream_payload && readStage_counterTwoValidStream_payload);
  assign when_SuperResolutionPart3_l500 = (readStage_counterTwoPixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart3_l502 = (readStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l504 = (readStage_mainThreeValidStream_payload && readStage_counterThreeValidStream_payload);
  assign when_SuperResolutionPart3_l511 = (readStage_counterThreePixelStream_payload <= readStage_mainThreePixelStream_payload);
  assign when_SuperResolutionPart3_l519 = (readStage_mainThreeValidStream_payload && readStage_counterOneValidStream_payload);
  assign when_SuperResolutionPart3_l521 = (readStage_mainOneValidStream_payload && readStage_counterThreeValidStream_payload);
  assign when_SuperResolutionPart3_l524 = (readStage_counterOnePixelStream_payload <= readStage_mainThreePixelStream_payload);
  assign when_SuperResolutionPart3_l526 = (readStage_counterThreePixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart3_l531 = (readStage_mainOneValidStream_payload && readStage_counterOneValidStream_payload);
  assign when_SuperResolutionPart3_l539 = (readStage_counterOnePixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart3_l547 = (readStage_mainOneValidStream_payload && readStage_counterThreeValidStream_payload);
  assign when_SuperResolutionPart3_l549 = (readStage_mainThreeValidStream_payload && readStage_counterOneValidStream_payload);
  assign when_SuperResolutionPart3_l552 = (readStage_counterThreePixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart3_l554 = (readStage_counterOnePixelStream_payload <= readStage_mainThreePixelStream_payload);
  assign when_SuperResolutionPart3_l559 = (readStage_mainThreeValidStream_payload && readStage_counterThreeValidStream_payload);
  assign when_SuperResolutionPart3_l562 = (readStage_counterThreePixelStream_payload <= readStage_mainThreePixelStream_payload);
  assign when_SuperResolutionPart3_l564 = (readStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l566 = (readStage_mainTwoValidStream_payload && readStage_counterTwoValidStream_payload);
  assign when_SuperResolutionPart3_l573 = (readStage_counterTwoPixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart3_l581 = (readStage_mainTwoValidStream_payload && readStage_counterOneValidStream_payload);
  assign when_SuperResolutionPart3_l583 = (readStage_mainOneValidStream_payload && readStage_counterTwoValidStream_payload);
  assign when_SuperResolutionPart3_l586 = (readStage_counterOnePixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart3_l588 = (readStage_counterTwoPixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart3_l593 = (readStage_mainOneValidStream_payload && readStage_counterOneValidStream_payload);
  assign when_SuperResolutionPart3_l601 = (readStage_counterOnePixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart3_l609 = (readStage_mainOneValidStream_payload && readStage_counterTwoValidStream_payload);
  assign when_SuperResolutionPart3_l611 = (readStage_mainTwoValidStream_payload && readStage_counterOneValidStream_payload);
  assign when_SuperResolutionPart3_l614 = (readStage_counterTwoPixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart3_l616 = (readStage_counterOnePixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart3_l496 = (readStage_controlPipe_payload_currentPosition == 2'b01);
  assign readStage_controlPipe_translated_valid = readStage_controlPipe_valid;
  assign readStage_controlPipe_ready = readStage_controlPipe_translated_ready;
  assign readStage_controlPipe_translated_payload_frameStart = readStage_controlPipe_payload_frameStart;
  assign readStage_controlPipe_translated_payload_rowEnd = readStage_controlPipe_payload_rowEnd;
  assign readStage_controlPipe_translated_payload_pipeValid = readStage_controlPipe_payload_pipeValid;
  assign readStage_controlPipe_translated_payload_firstRow = readStage_controlPipe_payload_firstRow;
  assign readStage_controlPipe_translated_payload_lastRow = readStage_controlPipe_payload_lastRow;
  assign readStage_controlPipe_translated_payload_finalResult = readStage_controlPipe_payload_finalResult;
  assign readStage_controlPipe_translated_payload_mainCompare = CICC1851_readStage_controlPipe_translated_payload_mainCompare;
  assign readStage_controlPipe_translated_payload_counterCompare = CICC1851_readStage_controlPipe_translated_payload_counterCompare;
  assign readStage_controlPipe_translated_payload_horizontalCompare = CICC1851_readStage_controlPipe_translated_payload_horizontalCompare;
  assign readStage_controlPipe_translated_payload_verticalCompare = CICC1851_readStage_controlPipe_translated_payload_verticalCompare;
  assign readStage_controlPipe_translated_payload_mainDiff = readStage_controlPipe_payload_mainDiff;
  assign readStage_controlPipe_translated_payload_counterDiff = readStage_controlPipe_payload_counterDiff;
  assign readStage_controlPipe_translated_payload_horizontalDiff = readStage_controlPipe_payload_horizontalDiff;
  assign readStage_controlPipe_translated_payload_verticalDiff = readStage_controlPipe_payload_verticalDiff;
  assign readStage_controlPipe_translated_payload_isHorizontalMin = readStage_controlPipe_payload_isHorizontalMin;
  assign readStage_controlPipe_translated_payload_minDiff = readStage_controlPipe_payload_minDiff;
  assign readStage_controlPipe_translated_payload_currentPosition = readStage_controlPipe_payload_currentPosition;
  assign readStage_controlPipe_translated_payload_nextPosition = readStage_controlPipe_payload_nextPosition;
  assign readStage_controlPipe_translated_payload_horizontalDirectionValid = CICC1851_readStage_controlPipe_translated_payload_horizontalDirectionValid;
  assign readStage_controlPipe_translated_payload_verticalDirectionValid = CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid;
  assign readStage_controlPipe_translated_payload_mainDirectionValid = CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid;
  assign readStage_controlPipe_translated_payload_counterDirectionValid = CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid;
  assign readStage_controlPipe_translated_payload_inValidMinDiff = readStage_controlPipe_payload_inValidMinDiff;
  assign readStage_controlPipe_translated_ready = (! readStage_controlPipe_translated_rValid);
  assign readStage_controlPipe_translated_s2mPipe_valid = (readStage_controlPipe_translated_valid || readStage_controlPipe_translated_rValid);
  assign readStage_controlPipe_translated_s2mPipe_payload_frameStart = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_frameStart : readStage_controlPipe_translated_payload_frameStart);
  assign readStage_controlPipe_translated_s2mPipe_payload_rowEnd = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_rowEnd : readStage_controlPipe_translated_payload_rowEnd);
  assign readStage_controlPipe_translated_s2mPipe_payload_pipeValid = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_pipeValid : readStage_controlPipe_translated_payload_pipeValid);
  assign readStage_controlPipe_translated_s2mPipe_payload_firstRow = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_firstRow : readStage_controlPipe_translated_payload_firstRow);
  assign readStage_controlPipe_translated_s2mPipe_payload_lastRow = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_lastRow : readStage_controlPipe_translated_payload_lastRow);
  assign readStage_controlPipe_translated_s2mPipe_payload_finalResult = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_finalResult : readStage_controlPipe_translated_payload_finalResult);
  assign readStage_controlPipe_translated_s2mPipe_payload_mainCompare = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_mainCompare : readStage_controlPipe_translated_payload_mainCompare);
  assign readStage_controlPipe_translated_s2mPipe_payload_counterCompare = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_counterCompare : readStage_controlPipe_translated_payload_counterCompare);
  assign readStage_controlPipe_translated_s2mPipe_payload_horizontalCompare = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_horizontalCompare : readStage_controlPipe_translated_payload_horizontalCompare);
  assign readStage_controlPipe_translated_s2mPipe_payload_verticalCompare = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_verticalCompare : readStage_controlPipe_translated_payload_verticalCompare);
  assign readStage_controlPipe_translated_s2mPipe_payload_mainDiff = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_mainDiff : readStage_controlPipe_translated_payload_mainDiff);
  assign readStage_controlPipe_translated_s2mPipe_payload_counterDiff = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_counterDiff : readStage_controlPipe_translated_payload_counterDiff);
  assign readStage_controlPipe_translated_s2mPipe_payload_horizontalDiff = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_horizontalDiff : readStage_controlPipe_translated_payload_horizontalDiff);
  assign readStage_controlPipe_translated_s2mPipe_payload_verticalDiff = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_verticalDiff : readStage_controlPipe_translated_payload_verticalDiff);
  assign readStage_controlPipe_translated_s2mPipe_payload_isHorizontalMin = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_isHorizontalMin : readStage_controlPipe_translated_payload_isHorizontalMin);
  assign readStage_controlPipe_translated_s2mPipe_payload_minDiff = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_minDiff : readStage_controlPipe_translated_payload_minDiff);
  assign readStage_controlPipe_translated_s2mPipe_payload_currentPosition = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_currentPosition : readStage_controlPipe_translated_payload_currentPosition);
  assign readStage_controlPipe_translated_s2mPipe_payload_nextPosition = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_nextPosition : readStage_controlPipe_translated_payload_nextPosition);
  assign readStage_controlPipe_translated_s2mPipe_payload_horizontalDirectionValid = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_horizontalDirectionValid : readStage_controlPipe_translated_payload_horizontalDirectionValid);
  assign readStage_controlPipe_translated_s2mPipe_payload_verticalDirectionValid = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_verticalDirectionValid : readStage_controlPipe_translated_payload_verticalDirectionValid);
  assign readStage_controlPipe_translated_s2mPipe_payload_mainDirectionValid = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_mainDirectionValid : readStage_controlPipe_translated_payload_mainDirectionValid);
  assign readStage_controlPipe_translated_s2mPipe_payload_counterDirectionValid = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_counterDirectionValid : readStage_controlPipe_translated_payload_counterDirectionValid);
  assign readStage_controlPipe_translated_s2mPipe_payload_inValidMinDiff = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_inValidMinDiff : readStage_controlPipe_translated_payload_inValidMinDiff);
  always @(*) begin
    readStage_controlPipe_translated_s2mPipe_ready = compareStage_controlPipe_ready;
    if(when_Stream_l368_40) begin
      readStage_controlPipe_translated_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_40 = (! compareStage_controlPipe_valid);
  assign compareStage_controlPipe_valid = readStage_controlPipe_translated_s2mPipe_rValid;
  assign compareStage_controlPipe_payload_frameStart = readStage_controlPipe_translated_s2mPipe_rData_frameStart;
  assign compareStage_controlPipe_payload_rowEnd = readStage_controlPipe_translated_s2mPipe_rData_rowEnd;
  assign compareStage_controlPipe_payload_pipeValid = readStage_controlPipe_translated_s2mPipe_rData_pipeValid;
  assign compareStage_controlPipe_payload_firstRow = readStage_controlPipe_translated_s2mPipe_rData_firstRow;
  assign compareStage_controlPipe_payload_lastRow = readStage_controlPipe_translated_s2mPipe_rData_lastRow;
  assign compareStage_controlPipe_payload_finalResult = readStage_controlPipe_translated_s2mPipe_rData_finalResult;
  assign compareStage_controlPipe_payload_mainCompare = readStage_controlPipe_translated_s2mPipe_rData_mainCompare;
  assign compareStage_controlPipe_payload_counterCompare = readStage_controlPipe_translated_s2mPipe_rData_counterCompare;
  assign compareStage_controlPipe_payload_horizontalCompare = readStage_controlPipe_translated_s2mPipe_rData_horizontalCompare;
  assign compareStage_controlPipe_payload_verticalCompare = readStage_controlPipe_translated_s2mPipe_rData_verticalCompare;
  assign compareStage_controlPipe_payload_mainDiff = readStage_controlPipe_translated_s2mPipe_rData_mainDiff;
  assign compareStage_controlPipe_payload_counterDiff = readStage_controlPipe_translated_s2mPipe_rData_counterDiff;
  assign compareStage_controlPipe_payload_horizontalDiff = readStage_controlPipe_translated_s2mPipe_rData_horizontalDiff;
  assign compareStage_controlPipe_payload_verticalDiff = readStage_controlPipe_translated_s2mPipe_rData_verticalDiff;
  assign compareStage_controlPipe_payload_isHorizontalMin = readStage_controlPipe_translated_s2mPipe_rData_isHorizontalMin;
  assign compareStage_controlPipe_payload_minDiff = readStage_controlPipe_translated_s2mPipe_rData_minDiff;
  assign compareStage_controlPipe_payload_currentPosition = readStage_controlPipe_translated_s2mPipe_rData_currentPosition;
  assign compareStage_controlPipe_payload_nextPosition = readStage_controlPipe_translated_s2mPipe_rData_nextPosition;
  assign compareStage_controlPipe_payload_horizontalDirectionValid = readStage_controlPipe_translated_s2mPipe_rData_horizontalDirectionValid;
  assign compareStage_controlPipe_payload_verticalDirectionValid = readStage_controlPipe_translated_s2mPipe_rData_verticalDirectionValid;
  assign compareStage_controlPipe_payload_mainDirectionValid = readStage_controlPipe_translated_s2mPipe_rData_mainDirectionValid;
  assign compareStage_controlPipe_payload_counterDirectionValid = readStage_controlPipe_translated_s2mPipe_rData_counterDirectionValid;
  assign compareStage_controlPipe_payload_inValidMinDiff = readStage_controlPipe_translated_s2mPipe_rData_inValidMinDiff;
  assign compareStage_mainOnePixelStream_ready = (! compareStage_mainOnePixelStream_rValid);
  assign compareStage_mainOnePixelStream_s2mPipe_valid = (compareStage_mainOnePixelStream_valid || compareStage_mainOnePixelStream_rValid);
  assign compareStage_mainOnePixelStream_s2mPipe_payload = (compareStage_mainOnePixelStream_rValid ? compareStage_mainOnePixelStream_rData : compareStage_mainOnePixelStream_payload);
  always @(*) begin
    compareStage_mainOnePixelStream_s2mPipe_ready = diffStage_mainOnePixelStream_ready;
    if(when_Stream_l368_41) begin
      compareStage_mainOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_41 = (! diffStage_mainOnePixelStream_valid);
  assign diffStage_mainOnePixelStream_valid = compareStage_mainOnePixelStream_s2mPipe_rValid;
  assign diffStage_mainOnePixelStream_payload = compareStage_mainOnePixelStream_s2mPipe_rData;
  assign compareStage_counterOnePixelStream_ready = (! compareStage_counterOnePixelStream_rValid);
  assign compareStage_counterOnePixelStream_s2mPipe_valid = (compareStage_counterOnePixelStream_valid || compareStage_counterOnePixelStream_rValid);
  assign compareStage_counterOnePixelStream_s2mPipe_payload = (compareStage_counterOnePixelStream_rValid ? compareStage_counterOnePixelStream_rData : compareStage_counterOnePixelStream_payload);
  always @(*) begin
    compareStage_counterOnePixelStream_s2mPipe_ready = diffStage_counterOnePixelStream_ready;
    if(when_Stream_l368_42) begin
      compareStage_counterOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_42 = (! diffStage_counterOnePixelStream_valid);
  assign diffStage_counterOnePixelStream_valid = compareStage_counterOnePixelStream_s2mPipe_rValid;
  assign diffStage_counterOnePixelStream_payload = compareStage_counterOnePixelStream_s2mPipe_rData;
  assign compareStage_mainTwoPixelStream_ready = (! compareStage_mainTwoPixelStream_rValid);
  assign compareStage_mainTwoPixelStream_s2mPipe_valid = (compareStage_mainTwoPixelStream_valid || compareStage_mainTwoPixelStream_rValid);
  assign compareStage_mainTwoPixelStream_s2mPipe_payload = (compareStage_mainTwoPixelStream_rValid ? compareStage_mainTwoPixelStream_rData : compareStage_mainTwoPixelStream_payload);
  always @(*) begin
    compareStage_mainTwoPixelStream_s2mPipe_ready = diffStage_mainTwoPixelStream_ready;
    if(when_Stream_l368_43) begin
      compareStage_mainTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_43 = (! diffStage_mainTwoPixelStream_valid);
  assign diffStage_mainTwoPixelStream_valid = compareStage_mainTwoPixelStream_s2mPipe_rValid;
  assign diffStage_mainTwoPixelStream_payload = compareStage_mainTwoPixelStream_s2mPipe_rData;
  assign compareStage_counterTwoPixelStream_ready = (! compareStage_counterTwoPixelStream_rValid);
  assign compareStage_counterTwoPixelStream_s2mPipe_valid = (compareStage_counterTwoPixelStream_valid || compareStage_counterTwoPixelStream_rValid);
  assign compareStage_counterTwoPixelStream_s2mPipe_payload = (compareStage_counterTwoPixelStream_rValid ? compareStage_counterTwoPixelStream_rData : compareStage_counterTwoPixelStream_payload);
  always @(*) begin
    compareStage_counterTwoPixelStream_s2mPipe_ready = diffStage_counterTwoPixelStream_ready;
    if(when_Stream_l368_44) begin
      compareStage_counterTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_44 = (! diffStage_counterTwoPixelStream_valid);
  assign diffStage_counterTwoPixelStream_valid = compareStage_counterTwoPixelStream_s2mPipe_rValid;
  assign diffStage_counterTwoPixelStream_payload = compareStage_counterTwoPixelStream_s2mPipe_rData;
  assign compareStage_mainThreePixelStream_ready = (! compareStage_mainThreePixelStream_rValid);
  assign compareStage_mainThreePixelStream_s2mPipe_valid = (compareStage_mainThreePixelStream_valid || compareStage_mainThreePixelStream_rValid);
  assign compareStage_mainThreePixelStream_s2mPipe_payload = (compareStage_mainThreePixelStream_rValid ? compareStage_mainThreePixelStream_rData : compareStage_mainThreePixelStream_payload);
  always @(*) begin
    compareStage_mainThreePixelStream_s2mPipe_ready = diffStage_mainThreePixelStream_ready;
    if(when_Stream_l368_45) begin
      compareStage_mainThreePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_45 = (! diffStage_mainThreePixelStream_valid);
  assign diffStage_mainThreePixelStream_valid = compareStage_mainThreePixelStream_s2mPipe_rValid;
  assign diffStage_mainThreePixelStream_payload = compareStage_mainThreePixelStream_s2mPipe_rData;
  assign compareStage_counterThreePixelStream_ready = (! compareStage_counterThreePixelStream_rValid);
  assign compareStage_counterThreePixelStream_s2mPipe_valid = (compareStage_counterThreePixelStream_valid || compareStage_counterThreePixelStream_rValid);
  assign compareStage_counterThreePixelStream_s2mPipe_payload = (compareStage_counterThreePixelStream_rValid ? compareStage_counterThreePixelStream_rData : compareStage_counterThreePixelStream_payload);
  always @(*) begin
    compareStage_counterThreePixelStream_s2mPipe_ready = diffStage_counterThreePixelStream_ready;
    if(when_Stream_l368_46) begin
      compareStage_counterThreePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_46 = (! diffStage_counterThreePixelStream_valid);
  assign diffStage_counterThreePixelStream_valid = compareStage_counterThreePixelStream_s2mPipe_rValid;
  assign diffStage_counterThreePixelStream_payload = compareStage_counterThreePixelStream_s2mPipe_rData;
  assign compareStage_mainOneValidStream_ready = (! compareStage_mainOneValidStream_rValid);
  assign compareStage_mainOneValidStream_s2mPipe_valid = (compareStage_mainOneValidStream_valid || compareStage_mainOneValidStream_rValid);
  assign compareStage_mainOneValidStream_s2mPipe_payload = (compareStage_mainOneValidStream_rValid ? compareStage_mainOneValidStream_rData : compareStage_mainOneValidStream_payload);
  always @(*) begin
    compareStage_mainOneValidStream_s2mPipe_ready = diffStage_mainOneValidStream_ready;
    if(when_Stream_l368_47) begin
      compareStage_mainOneValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_47 = (! diffStage_mainOneValidStream_valid);
  assign diffStage_mainOneValidStream_valid = compareStage_mainOneValidStream_s2mPipe_rValid;
  assign diffStage_mainOneValidStream_payload = compareStage_mainOneValidStream_s2mPipe_rData;
  assign compareStage_counterOneValidStream_ready = (! compareStage_counterOneValidStream_rValid);
  assign compareStage_counterOneValidStream_s2mPipe_valid = (compareStage_counterOneValidStream_valid || compareStage_counterOneValidStream_rValid);
  assign compareStage_counterOneValidStream_s2mPipe_payload = (compareStage_counterOneValidStream_rValid ? compareStage_counterOneValidStream_rData : compareStage_counterOneValidStream_payload);
  always @(*) begin
    compareStage_counterOneValidStream_s2mPipe_ready = diffStage_counterOneValidStream_ready;
    if(when_Stream_l368_48) begin
      compareStage_counterOneValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_48 = (! diffStage_counterOneValidStream_valid);
  assign diffStage_counterOneValidStream_valid = compareStage_counterOneValidStream_s2mPipe_rValid;
  assign diffStage_counterOneValidStream_payload = compareStage_counterOneValidStream_s2mPipe_rData;
  assign compareStage_mainTwoValidStream_ready = (! compareStage_mainTwoValidStream_rValid);
  assign compareStage_mainTwoValidStream_s2mPipe_valid = (compareStage_mainTwoValidStream_valid || compareStage_mainTwoValidStream_rValid);
  assign compareStage_mainTwoValidStream_s2mPipe_payload = (compareStage_mainTwoValidStream_rValid ? compareStage_mainTwoValidStream_rData : compareStage_mainTwoValidStream_payload);
  always @(*) begin
    compareStage_mainTwoValidStream_s2mPipe_ready = diffStage_mainTwoValidStream_ready;
    if(when_Stream_l368_49) begin
      compareStage_mainTwoValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_49 = (! diffStage_mainTwoValidStream_valid);
  assign diffStage_mainTwoValidStream_valid = compareStage_mainTwoValidStream_s2mPipe_rValid;
  assign diffStage_mainTwoValidStream_payload = compareStage_mainTwoValidStream_s2mPipe_rData;
  assign compareStage_counterTwoValidStream_ready = (! compareStage_counterTwoValidStream_rValid);
  assign compareStage_counterTwoValidStream_s2mPipe_valid = (compareStage_counterTwoValidStream_valid || compareStage_counterTwoValidStream_rValid);
  assign compareStage_counterTwoValidStream_s2mPipe_payload = (compareStage_counterTwoValidStream_rValid ? compareStage_counterTwoValidStream_rData : compareStage_counterTwoValidStream_payload);
  always @(*) begin
    compareStage_counterTwoValidStream_s2mPipe_ready = diffStage_counterTwoValidStream_ready;
    if(when_Stream_l368_50) begin
      compareStage_counterTwoValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_50 = (! diffStage_counterTwoValidStream_valid);
  assign diffStage_counterTwoValidStream_valid = compareStage_counterTwoValidStream_s2mPipe_rValid;
  assign diffStage_counterTwoValidStream_payload = compareStage_counterTwoValidStream_s2mPipe_rData;
  assign compareStage_mainThreeValidStream_ready = (! compareStage_mainThreeValidStream_rValid);
  assign compareStage_mainThreeValidStream_s2mPipe_valid = (compareStage_mainThreeValidStream_valid || compareStage_mainThreeValidStream_rValid);
  assign compareStage_mainThreeValidStream_s2mPipe_payload = (compareStage_mainThreeValidStream_rValid ? compareStage_mainThreeValidStream_rData : compareStage_mainThreeValidStream_payload);
  always @(*) begin
    compareStage_mainThreeValidStream_s2mPipe_ready = diffStage_mainThreeValidStream_ready;
    if(when_Stream_l368_51) begin
      compareStage_mainThreeValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_51 = (! diffStage_mainThreeValidStream_valid);
  assign diffStage_mainThreeValidStream_valid = compareStage_mainThreeValidStream_s2mPipe_rValid;
  assign diffStage_mainThreeValidStream_payload = compareStage_mainThreeValidStream_s2mPipe_rData;
  assign compareStage_counterThreeValidStream_ready = (! compareStage_counterThreeValidStream_rValid);
  assign compareStage_counterThreeValidStream_s2mPipe_valid = (compareStage_counterThreeValidStream_valid || compareStage_counterThreeValidStream_rValid);
  assign compareStage_counterThreeValidStream_s2mPipe_payload = (compareStage_counterThreeValidStream_rValid ? compareStage_counterThreeValidStream_rData : compareStage_counterThreeValidStream_payload);
  always @(*) begin
    compareStage_counterThreeValidStream_s2mPipe_ready = diffStage_counterThreeValidStream_ready;
    if(when_Stream_l368_52) begin
      compareStage_counterThreeValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_52 = (! diffStage_counterThreeValidStream_valid);
  assign diffStage_counterThreeValidStream_valid = compareStage_counterThreeValidStream_s2mPipe_rValid;
  assign diffStage_counterThreeValidStream_payload = compareStage_counterThreeValidStream_s2mPipe_rData;
  always @(*) begin
    CICC1851_compareStage_controlPipe_translated_payload_mainDiff = compareStage_controlPipe_payload_mainDiff;
    if(!compareStage_controlPipe_payload_finalResult) begin
      if(when_SuperResolutionPart3_l661) begin
        if(when_SuperResolutionPart3_l664) begin
          if(compareStage_controlPipe_payload_firstRow) begin
            if(compareStage_controlPipe_payload_mainCompare) begin
              CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterTwoPixelStream_payload);
            end else begin
              CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainTwoPixelStream_payload);
            end
          end else begin
            if(compareStage_controlPipe_payload_lastRow) begin
              if(compareStage_controlPipe_payload_mainCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainThreePixelStream_payload - compareStage_counterThreePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterThreePixelStream_payload - compareStage_mainThreePixelStream_payload);
              end
            end else begin
              if(compareStage_controlPipe_payload_mainCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainThreePixelStream_payload - compareStage_counterTwoPixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainThreePixelStream_payload);
              end
            end
          end
        end else begin
          if(compareStage_controlPipe_payload_lastRow) begin
            if(compareStage_controlPipe_payload_mainCompare) begin
              CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterTwoPixelStream_payload);
            end else begin
              CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainTwoPixelStream_payload);
            end
          end else begin
            if(compareStage_controlPipe_payload_mainCompare) begin
              CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterThreePixelStream_payload);
            end else begin
              CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterThreePixelStream_payload - compareStage_mainTwoPixelStream_payload);
            end
          end
        end
      end else begin
        if(when_SuperResolutionPart3_l694) begin
          if(when_SuperResolutionPart3_l697) begin
            if(compareStage_controlPipe_payload_lastRow) begin
              if(compareStage_controlPipe_payload_mainCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainThreePixelStream_payload - compareStage_counterThreePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterThreePixelStream_payload - compareStage_mainThreePixelStream_payload);
              end
            end else begin
              if(compareStage_controlPipe_payload_mainCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainThreePixelStream_payload - compareStage_counterOnePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterOnePixelStream_payload - compareStage_mainThreePixelStream_payload);
              end
            end
          end else begin
            if(compareStage_controlPipe_payload_lastRow) begin
              if(compareStage_controlPipe_payload_mainCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_counterOnePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterOnePixelStream_payload - compareStage_mainOnePixelStream_payload);
              end
            end else begin
              if(compareStage_controlPipe_payload_mainCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_counterThreePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterThreePixelStream_payload - compareStage_mainOnePixelStream_payload);
              end
            end
          end
        end else begin
          if(when_SuperResolutionPart3_l725) begin
            if(compareStage_controlPipe_payload_lastRow) begin
              if(compareStage_controlPipe_payload_mainCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterTwoPixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainTwoPixelStream_payload);
              end
            end else begin
              if(compareStage_controlPipe_payload_mainCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterOnePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterOnePixelStream_payload - compareStage_mainTwoPixelStream_payload);
              end
            end
          end else begin
            if(compareStage_controlPipe_payload_lastRow) begin
              if(compareStage_controlPipe_payload_mainCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_counterOnePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterOnePixelStream_payload - compareStage_mainOnePixelStream_payload);
              end
            end else begin
              if(compareStage_controlPipe_payload_mainCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_counterTwoPixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainOnePixelStream_payload);
              end
            end
          end
        end
      end
    end
  end

  always @(*) begin
    CICC1851_compareStage_controlPipe_translated_payload_counterDiff = compareStage_controlPipe_payload_counterDiff;
    if(!compareStage_controlPipe_payload_finalResult) begin
      if(when_SuperResolutionPart3_l661) begin
        if(when_SuperResolutionPart3_l664) begin
          if(compareStage_controlPipe_payload_firstRow) begin
            if(compareStage_controlPipe_payload_counterCompare) begin
              CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterTwoPixelStream_payload);
            end else begin
              CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainTwoPixelStream_payload);
            end
          end else begin
            if(compareStage_controlPipe_payload_lastRow) begin
              if(compareStage_controlPipe_payload_counterCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_mainThreePixelStream_payload - compareStage_counterThreePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterThreePixelStream_payload - compareStage_mainThreePixelStream_payload);
              end
            end else begin
              if(compareStage_controlPipe_payload_counterCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterThreePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterThreePixelStream_payload - compareStage_mainTwoPixelStream_payload);
              end
            end
          end
        end else begin
          if(compareStage_controlPipe_payload_lastRow) begin
            if(compareStage_controlPipe_payload_counterCompare) begin
              CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterTwoPixelStream_payload);
            end else begin
              CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainTwoPixelStream_payload);
            end
          end else begin
            if(compareStage_controlPipe_payload_counterCompare) begin
              CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_mainThreePixelStream_payload - compareStage_counterTwoPixelStream_payload);
            end else begin
              CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainThreePixelStream_payload);
            end
          end
        end
      end else begin
        if(when_SuperResolutionPart3_l694) begin
          if(when_SuperResolutionPart3_l697) begin
            if(compareStage_controlPipe_payload_lastRow) begin
              if(compareStage_controlPipe_payload_counterCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_mainThreePixelStream_payload - compareStage_counterThreePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterThreePixelStream_payload - compareStage_mainThreePixelStream_payload);
              end
            end else begin
              if(compareStage_controlPipe_payload_counterCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_mainOnePixelStream_payload - compareStage_counterThreePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterThreePixelStream_payload - compareStage_mainOnePixelStream_payload);
              end
            end
          end else begin
            if(compareStage_controlPipe_payload_lastRow) begin
              if(compareStage_controlPipe_payload_counterCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_mainOnePixelStream_payload - compareStage_counterOnePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterOnePixelStream_payload - compareStage_mainOnePixelStream_payload);
              end
            end else begin
              if(compareStage_controlPipe_payload_counterCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_mainThreePixelStream_payload - compareStage_counterOnePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterOnePixelStream_payload - compareStage_mainThreePixelStream_payload);
              end
            end
          end
        end else begin
          if(when_SuperResolutionPart3_l725) begin
            if(compareStage_controlPipe_payload_lastRow) begin
              if(compareStage_controlPipe_payload_counterCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterTwoPixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainTwoPixelStream_payload);
              end
            end else begin
              if(compareStage_controlPipe_payload_counterCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_mainOnePixelStream_payload - compareStage_counterTwoPixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainOnePixelStream_payload);
              end
            end
          end else begin
            if(compareStage_controlPipe_payload_lastRow) begin
              if(compareStage_controlPipe_payload_counterCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_mainOnePixelStream_payload - compareStage_counterOnePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterOnePixelStream_payload - compareStage_mainOnePixelStream_payload);
              end
            end else begin
              if(compareStage_controlPipe_payload_counterCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterOnePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterOnePixelStream_payload - compareStage_mainTwoPixelStream_payload);
              end
            end
          end
        end
      end
    end
  end

  always @(*) begin
    CICC1851_compareStage_controlPipe_translated_payload_horizontalDiff = compareStage_controlPipe_payload_horizontalDiff;
    if(!compareStage_controlPipe_payload_finalResult) begin
      if(when_SuperResolutionPart3_l661) begin
        if(compareStage_controlPipe_payload_horizontalCompare) begin
          CICC1851_compareStage_controlPipe_translated_payload_horizontalDiff = (compareStage_mainOnePixelStream_payload - compareStage_counterOnePixelStream_payload);
        end else begin
          CICC1851_compareStage_controlPipe_translated_payload_horizontalDiff = (compareStage_counterOnePixelStream_payload - compareStage_mainOnePixelStream_payload);
        end
      end else begin
        if(when_SuperResolutionPart3_l694) begin
          if(compareStage_controlPipe_payload_horizontalCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_horizontalDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterTwoPixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_horizontalDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainTwoPixelStream_payload);
          end
        end else begin
          if(compareStage_controlPipe_payload_horizontalCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_horizontalDiff = (compareStage_mainThreePixelStream_payload - compareStage_counterThreePixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_horizontalDiff = (compareStage_counterThreePixelStream_payload - compareStage_mainThreePixelStream_payload);
          end
        end
      end
    end
  end

  always @(*) begin
    CICC1851_compareStage_controlPipe_translated_payload_verticalDiff = compareStage_controlPipe_payload_verticalDiff;
    if(compareStage_controlPipe_payload_finalResult) begin
      if(when_SuperResolutionPart3_l647) begin
        CICC1851_compareStage_controlPipe_translated_payload_verticalDiff = 8'h0;
      end else begin
        if(when_SuperResolutionPart3_l649) begin
          if(compareStage_controlPipe_payload_verticalCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_verticalDiff = (compareStage_mainTwoPixelStream_payload - compareStage_mainThreePixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_verticalDiff = (compareStage_mainThreePixelStream_payload - compareStage_mainTwoPixelStream_payload);
          end
        end else begin
          if(when_SuperResolutionPart3_l652) begin
            if(compareStage_controlPipe_payload_verticalCompare) begin
              CICC1851_compareStage_controlPipe_translated_payload_verticalDiff = (compareStage_mainOnePixelStream_payload - compareStage_mainThreePixelStream_payload);
            end else begin
              CICC1851_compareStage_controlPipe_translated_payload_verticalDiff = (compareStage_mainThreePixelStream_payload - compareStage_mainOnePixelStream_payload);
            end
          end else begin
            if(compareStage_controlPipe_payload_verticalCompare) begin
              CICC1851_compareStage_controlPipe_translated_payload_verticalDiff = (compareStage_mainOnePixelStream_payload - compareStage_mainTwoPixelStream_payload);
            end else begin
              CICC1851_compareStage_controlPipe_translated_payload_verticalDiff = (compareStage_mainTwoPixelStream_payload - compareStage_mainOnePixelStream_payload);
            end
          end
        end
      end
    end
  end

  always @(*) begin
    CICC1851_compareStage_controlPipe_translated_payload_inValidMinDiff = compareStage_controlPipe_payload_inValidMinDiff;
    if(when_SuperResolutionPart3_l753) begin
      CICC1851_compareStage_controlPipe_translated_payload_inValidMinDiff = 1'b1;
    end
  end

  assign when_SuperResolutionPart3_l647 = (compareStage_controlPipe_payload_firstRow || compareStage_controlPipe_payload_lastRow);
  assign when_SuperResolutionPart3_l649 = (compareStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l652 = (compareStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l661 = (compareStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l664 = (compareStage_controlPipe_payload_nextPosition == 2'b01);
  assign when_SuperResolutionPart3_l697 = (compareStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l725 = (compareStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l694 = (compareStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l753 = ((((! compareStage_controlPipe_payload_finalResult) && (! compareStage_controlPipe_payload_mainDirectionValid)) && (! compareStage_controlPipe_payload_counterDirectionValid)) && (! compareStage_controlPipe_payload_horizontalDirectionValid));
  assign compareStage_controlPipe_translated_valid = compareStage_controlPipe_valid;
  assign compareStage_controlPipe_ready = compareStage_controlPipe_translated_ready;
  assign compareStage_controlPipe_translated_payload_frameStart = compareStage_controlPipe_payload_frameStart;
  assign compareStage_controlPipe_translated_payload_rowEnd = compareStage_controlPipe_payload_rowEnd;
  assign compareStage_controlPipe_translated_payload_pipeValid = compareStage_controlPipe_payload_pipeValid;
  assign compareStage_controlPipe_translated_payload_firstRow = compareStage_controlPipe_payload_firstRow;
  assign compareStage_controlPipe_translated_payload_lastRow = compareStage_controlPipe_payload_lastRow;
  assign compareStage_controlPipe_translated_payload_finalResult = compareStage_controlPipe_payload_finalResult;
  assign compareStage_controlPipe_translated_payload_mainCompare = compareStage_controlPipe_payload_mainCompare;
  assign compareStage_controlPipe_translated_payload_counterCompare = compareStage_controlPipe_payload_counterCompare;
  assign compareStage_controlPipe_translated_payload_horizontalCompare = compareStage_controlPipe_payload_horizontalCompare;
  assign compareStage_controlPipe_translated_payload_verticalCompare = compareStage_controlPipe_payload_verticalCompare;
  assign compareStage_controlPipe_translated_payload_mainDiff = CICC1851_compareStage_controlPipe_translated_payload_mainDiff;
  assign compareStage_controlPipe_translated_payload_counterDiff = CICC1851_compareStage_controlPipe_translated_payload_counterDiff;
  assign compareStage_controlPipe_translated_payload_horizontalDiff = CICC1851_compareStage_controlPipe_translated_payload_horizontalDiff;
  assign compareStage_controlPipe_translated_payload_verticalDiff = CICC1851_compareStage_controlPipe_translated_payload_verticalDiff;
  assign compareStage_controlPipe_translated_payload_isHorizontalMin = compareStage_controlPipe_payload_isHorizontalMin;
  assign compareStage_controlPipe_translated_payload_minDiff = compareStage_controlPipe_payload_minDiff;
  assign compareStage_controlPipe_translated_payload_currentPosition = compareStage_controlPipe_payload_currentPosition;
  assign compareStage_controlPipe_translated_payload_nextPosition = compareStage_controlPipe_payload_nextPosition;
  assign compareStage_controlPipe_translated_payload_horizontalDirectionValid = compareStage_controlPipe_payload_horizontalDirectionValid;
  assign compareStage_controlPipe_translated_payload_verticalDirectionValid = compareStage_controlPipe_payload_verticalDirectionValid;
  assign compareStage_controlPipe_translated_payload_mainDirectionValid = compareStage_controlPipe_payload_mainDirectionValid;
  assign compareStage_controlPipe_translated_payload_counterDirectionValid = compareStage_controlPipe_payload_counterDirectionValid;
  assign compareStage_controlPipe_translated_payload_inValidMinDiff = CICC1851_compareStage_controlPipe_translated_payload_inValidMinDiff;
  assign compareStage_controlPipe_translated_ready = (! compareStage_controlPipe_translated_rValid);
  assign compareStage_controlPipe_translated_s2mPipe_valid = (compareStage_controlPipe_translated_valid || compareStage_controlPipe_translated_rValid);
  assign compareStage_controlPipe_translated_s2mPipe_payload_frameStart = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_frameStart : compareStage_controlPipe_translated_payload_frameStart);
  assign compareStage_controlPipe_translated_s2mPipe_payload_rowEnd = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_rowEnd : compareStage_controlPipe_translated_payload_rowEnd);
  assign compareStage_controlPipe_translated_s2mPipe_payload_pipeValid = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_pipeValid : compareStage_controlPipe_translated_payload_pipeValid);
  assign compareStage_controlPipe_translated_s2mPipe_payload_firstRow = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_firstRow : compareStage_controlPipe_translated_payload_firstRow);
  assign compareStage_controlPipe_translated_s2mPipe_payload_lastRow = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_lastRow : compareStage_controlPipe_translated_payload_lastRow);
  assign compareStage_controlPipe_translated_s2mPipe_payload_finalResult = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_finalResult : compareStage_controlPipe_translated_payload_finalResult);
  assign compareStage_controlPipe_translated_s2mPipe_payload_mainCompare = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_mainCompare : compareStage_controlPipe_translated_payload_mainCompare);
  assign compareStage_controlPipe_translated_s2mPipe_payload_counterCompare = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_counterCompare : compareStage_controlPipe_translated_payload_counterCompare);
  assign compareStage_controlPipe_translated_s2mPipe_payload_horizontalCompare = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_horizontalCompare : compareStage_controlPipe_translated_payload_horizontalCompare);
  assign compareStage_controlPipe_translated_s2mPipe_payload_verticalCompare = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_verticalCompare : compareStage_controlPipe_translated_payload_verticalCompare);
  assign compareStage_controlPipe_translated_s2mPipe_payload_mainDiff = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_mainDiff : compareStage_controlPipe_translated_payload_mainDiff);
  assign compareStage_controlPipe_translated_s2mPipe_payload_counterDiff = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_counterDiff : compareStage_controlPipe_translated_payload_counterDiff);
  assign compareStage_controlPipe_translated_s2mPipe_payload_horizontalDiff = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_horizontalDiff : compareStage_controlPipe_translated_payload_horizontalDiff);
  assign compareStage_controlPipe_translated_s2mPipe_payload_verticalDiff = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_verticalDiff : compareStage_controlPipe_translated_payload_verticalDiff);
  assign compareStage_controlPipe_translated_s2mPipe_payload_isHorizontalMin = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_isHorizontalMin : compareStage_controlPipe_translated_payload_isHorizontalMin);
  assign compareStage_controlPipe_translated_s2mPipe_payload_minDiff = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_minDiff : compareStage_controlPipe_translated_payload_minDiff);
  assign compareStage_controlPipe_translated_s2mPipe_payload_currentPosition = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_currentPosition : compareStage_controlPipe_translated_payload_currentPosition);
  assign compareStage_controlPipe_translated_s2mPipe_payload_nextPosition = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_nextPosition : compareStage_controlPipe_translated_payload_nextPosition);
  assign compareStage_controlPipe_translated_s2mPipe_payload_horizontalDirectionValid = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_horizontalDirectionValid : compareStage_controlPipe_translated_payload_horizontalDirectionValid);
  assign compareStage_controlPipe_translated_s2mPipe_payload_verticalDirectionValid = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_verticalDirectionValid : compareStage_controlPipe_translated_payload_verticalDirectionValid);
  assign compareStage_controlPipe_translated_s2mPipe_payload_mainDirectionValid = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_mainDirectionValid : compareStage_controlPipe_translated_payload_mainDirectionValid);
  assign compareStage_controlPipe_translated_s2mPipe_payload_counterDirectionValid = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_counterDirectionValid : compareStage_controlPipe_translated_payload_counterDirectionValid);
  assign compareStage_controlPipe_translated_s2mPipe_payload_inValidMinDiff = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_inValidMinDiff : compareStage_controlPipe_translated_payload_inValidMinDiff);
  always @(*) begin
    compareStage_controlPipe_translated_s2mPipe_ready = diffStage_controlPipe_ready;
    if(when_Stream_l368_53) begin
      compareStage_controlPipe_translated_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_53 = (! diffStage_controlPipe_valid);
  assign diffStage_controlPipe_valid = compareStage_controlPipe_translated_s2mPipe_rValid;
  assign diffStage_controlPipe_payload_frameStart = compareStage_controlPipe_translated_s2mPipe_rData_frameStart;
  assign diffStage_controlPipe_payload_rowEnd = compareStage_controlPipe_translated_s2mPipe_rData_rowEnd;
  assign diffStage_controlPipe_payload_pipeValid = compareStage_controlPipe_translated_s2mPipe_rData_pipeValid;
  assign diffStage_controlPipe_payload_firstRow = compareStage_controlPipe_translated_s2mPipe_rData_firstRow;
  assign diffStage_controlPipe_payload_lastRow = compareStage_controlPipe_translated_s2mPipe_rData_lastRow;
  assign diffStage_controlPipe_payload_finalResult = compareStage_controlPipe_translated_s2mPipe_rData_finalResult;
  assign diffStage_controlPipe_payload_mainCompare = compareStage_controlPipe_translated_s2mPipe_rData_mainCompare;
  assign diffStage_controlPipe_payload_counterCompare = compareStage_controlPipe_translated_s2mPipe_rData_counterCompare;
  assign diffStage_controlPipe_payload_horizontalCompare = compareStage_controlPipe_translated_s2mPipe_rData_horizontalCompare;
  assign diffStage_controlPipe_payload_verticalCompare = compareStage_controlPipe_translated_s2mPipe_rData_verticalCompare;
  assign diffStage_controlPipe_payload_mainDiff = compareStage_controlPipe_translated_s2mPipe_rData_mainDiff;
  assign diffStage_controlPipe_payload_counterDiff = compareStage_controlPipe_translated_s2mPipe_rData_counterDiff;
  assign diffStage_controlPipe_payload_horizontalDiff = compareStage_controlPipe_translated_s2mPipe_rData_horizontalDiff;
  assign diffStage_controlPipe_payload_verticalDiff = compareStage_controlPipe_translated_s2mPipe_rData_verticalDiff;
  assign diffStage_controlPipe_payload_isHorizontalMin = compareStage_controlPipe_translated_s2mPipe_rData_isHorizontalMin;
  assign diffStage_controlPipe_payload_minDiff = compareStage_controlPipe_translated_s2mPipe_rData_minDiff;
  assign diffStage_controlPipe_payload_currentPosition = compareStage_controlPipe_translated_s2mPipe_rData_currentPosition;
  assign diffStage_controlPipe_payload_nextPosition = compareStage_controlPipe_translated_s2mPipe_rData_nextPosition;
  assign diffStage_controlPipe_payload_horizontalDirectionValid = compareStage_controlPipe_translated_s2mPipe_rData_horizontalDirectionValid;
  assign diffStage_controlPipe_payload_verticalDirectionValid = compareStage_controlPipe_translated_s2mPipe_rData_verticalDirectionValid;
  assign diffStage_controlPipe_payload_mainDirectionValid = compareStage_controlPipe_translated_s2mPipe_rData_mainDirectionValid;
  assign diffStage_controlPipe_payload_counterDirectionValid = compareStage_controlPipe_translated_s2mPipe_rData_counterDirectionValid;
  assign diffStage_controlPipe_payload_inValidMinDiff = compareStage_controlPipe_translated_s2mPipe_rData_inValidMinDiff;
  assign diffStage_mainOnePixelStream_ready = (! diffStage_mainOnePixelStream_rValid);
  assign diffStage_mainOnePixelStream_s2mPipe_valid = (diffStage_mainOnePixelStream_valid || diffStage_mainOnePixelStream_rValid);
  assign diffStage_mainOnePixelStream_s2mPipe_payload = (diffStage_mainOnePixelStream_rValid ? diffStage_mainOnePixelStream_rData : diffStage_mainOnePixelStream_payload);
  always @(*) begin
    diffStage_mainOnePixelStream_s2mPipe_ready = resultStage_mainOnePixelStream_ready;
    if(when_Stream_l368_54) begin
      diffStage_mainOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_54 = (! resultStage_mainOnePixelStream_valid);
  assign resultStage_mainOnePixelStream_valid = diffStage_mainOnePixelStream_s2mPipe_rValid;
  assign resultStage_mainOnePixelStream_payload = diffStage_mainOnePixelStream_s2mPipe_rData;
  assign diffStage_counterOnePixelStream_ready = (! diffStage_counterOnePixelStream_rValid);
  assign diffStage_counterOnePixelStream_s2mPipe_valid = (diffStage_counterOnePixelStream_valid || diffStage_counterOnePixelStream_rValid);
  assign diffStage_counterOnePixelStream_s2mPipe_payload = (diffStage_counterOnePixelStream_rValid ? diffStage_counterOnePixelStream_rData : diffStage_counterOnePixelStream_payload);
  always @(*) begin
    diffStage_counterOnePixelStream_s2mPipe_ready = resultStage_counterOnePixelStream_ready;
    if(when_Stream_l368_55) begin
      diffStage_counterOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_55 = (! resultStage_counterOnePixelStream_valid);
  assign resultStage_counterOnePixelStream_valid = diffStage_counterOnePixelStream_s2mPipe_rValid;
  assign resultStage_counterOnePixelStream_payload = diffStage_counterOnePixelStream_s2mPipe_rData;
  assign diffStage_mainTwoPixelStream_ready = (! diffStage_mainTwoPixelStream_rValid);
  assign diffStage_mainTwoPixelStream_s2mPipe_valid = (diffStage_mainTwoPixelStream_valid || diffStage_mainTwoPixelStream_rValid);
  assign diffStage_mainTwoPixelStream_s2mPipe_payload = (diffStage_mainTwoPixelStream_rValid ? diffStage_mainTwoPixelStream_rData : diffStage_mainTwoPixelStream_payload);
  always @(*) begin
    diffStage_mainTwoPixelStream_s2mPipe_ready = resultStage_mainTwoPixelStream_ready;
    if(when_Stream_l368_56) begin
      diffStage_mainTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_56 = (! resultStage_mainTwoPixelStream_valid);
  assign resultStage_mainTwoPixelStream_valid = diffStage_mainTwoPixelStream_s2mPipe_rValid;
  assign resultStage_mainTwoPixelStream_payload = diffStage_mainTwoPixelStream_s2mPipe_rData;
  assign diffStage_counterTwoPixelStream_ready = (! diffStage_counterTwoPixelStream_rValid);
  assign diffStage_counterTwoPixelStream_s2mPipe_valid = (diffStage_counterTwoPixelStream_valid || diffStage_counterTwoPixelStream_rValid);
  assign diffStage_counterTwoPixelStream_s2mPipe_payload = (diffStage_counterTwoPixelStream_rValid ? diffStage_counterTwoPixelStream_rData : diffStage_counterTwoPixelStream_payload);
  always @(*) begin
    diffStage_counterTwoPixelStream_s2mPipe_ready = resultStage_counterTwoPixelStream_ready;
    if(when_Stream_l368_57) begin
      diffStage_counterTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_57 = (! resultStage_counterTwoPixelStream_valid);
  assign resultStage_counterTwoPixelStream_valid = diffStage_counterTwoPixelStream_s2mPipe_rValid;
  assign resultStage_counterTwoPixelStream_payload = diffStage_counterTwoPixelStream_s2mPipe_rData;
  assign diffStage_mainThreePixelStream_ready = (! diffStage_mainThreePixelStream_rValid);
  assign diffStage_mainThreePixelStream_s2mPipe_valid = (diffStage_mainThreePixelStream_valid || diffStage_mainThreePixelStream_rValid);
  assign diffStage_mainThreePixelStream_s2mPipe_payload = (diffStage_mainThreePixelStream_rValid ? diffStage_mainThreePixelStream_rData : diffStage_mainThreePixelStream_payload);
  always @(*) begin
    diffStage_mainThreePixelStream_s2mPipe_ready = resultStage_mainThreePixelStream_ready;
    if(when_Stream_l368_58) begin
      diffStage_mainThreePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_58 = (! resultStage_mainThreePixelStream_valid);
  assign resultStage_mainThreePixelStream_valid = diffStage_mainThreePixelStream_s2mPipe_rValid;
  assign resultStage_mainThreePixelStream_payload = diffStage_mainThreePixelStream_s2mPipe_rData;
  assign diffStage_counterThreePixelStream_ready = (! diffStage_counterThreePixelStream_rValid);
  assign diffStage_counterThreePixelStream_s2mPipe_valid = (diffStage_counterThreePixelStream_valid || diffStage_counterThreePixelStream_rValid);
  assign diffStage_counterThreePixelStream_s2mPipe_payload = (diffStage_counterThreePixelStream_rValid ? diffStage_counterThreePixelStream_rData : diffStage_counterThreePixelStream_payload);
  always @(*) begin
    diffStage_counterThreePixelStream_s2mPipe_ready = resultStage_counterThreePixelStream_ready;
    if(when_Stream_l368_59) begin
      diffStage_counterThreePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_59 = (! resultStage_counterThreePixelStream_valid);
  assign resultStage_counterThreePixelStream_valid = diffStage_counterThreePixelStream_s2mPipe_rValid;
  assign resultStage_counterThreePixelStream_payload = diffStage_counterThreePixelStream_s2mPipe_rData;
  assign diffStage_mainOneValidStream_ready = (! diffStage_mainOneValidStream_rValid);
  assign diffStage_mainOneValidStream_s2mPipe_valid = (diffStage_mainOneValidStream_valid || diffStage_mainOneValidStream_rValid);
  assign diffStage_mainOneValidStream_s2mPipe_payload = (diffStage_mainOneValidStream_rValid ? diffStage_mainOneValidStream_rData : diffStage_mainOneValidStream_payload);
  always @(*) begin
    diffStage_mainOneValidStream_s2mPipe_ready = resultStage_mainOneValidStream_ready;
    if(when_Stream_l368_60) begin
      diffStage_mainOneValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_60 = (! resultStage_mainOneValidStream_valid);
  assign resultStage_mainOneValidStream_valid = diffStage_mainOneValidStream_s2mPipe_rValid;
  assign resultStage_mainOneValidStream_payload = diffStage_mainOneValidStream_s2mPipe_rData;
  assign diffStage_counterOneValidStream_ready = (! diffStage_counterOneValidStream_rValid);
  assign diffStage_counterOneValidStream_s2mPipe_valid = (diffStage_counterOneValidStream_valid || diffStage_counterOneValidStream_rValid);
  assign diffStage_counterOneValidStream_s2mPipe_payload = (diffStage_counterOneValidStream_rValid ? diffStage_counterOneValidStream_rData : diffStage_counterOneValidStream_payload);
  always @(*) begin
    diffStage_counterOneValidStream_s2mPipe_ready = resultStage_counterOneValidStream_ready;
    if(when_Stream_l368_61) begin
      diffStage_counterOneValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_61 = (! resultStage_counterOneValidStream_valid);
  assign resultStage_counterOneValidStream_valid = diffStage_counterOneValidStream_s2mPipe_rValid;
  assign resultStage_counterOneValidStream_payload = diffStage_counterOneValidStream_s2mPipe_rData;
  assign diffStage_mainTwoValidStream_ready = (! diffStage_mainTwoValidStream_rValid);
  assign diffStage_mainTwoValidStream_s2mPipe_valid = (diffStage_mainTwoValidStream_valid || diffStage_mainTwoValidStream_rValid);
  assign diffStage_mainTwoValidStream_s2mPipe_payload = (diffStage_mainTwoValidStream_rValid ? diffStage_mainTwoValidStream_rData : diffStage_mainTwoValidStream_payload);
  always @(*) begin
    diffStage_mainTwoValidStream_s2mPipe_ready = resultStage_mainTwoValidStream_ready;
    if(when_Stream_l368_62) begin
      diffStage_mainTwoValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_62 = (! resultStage_mainTwoValidStream_valid);
  assign resultStage_mainTwoValidStream_valid = diffStage_mainTwoValidStream_s2mPipe_rValid;
  assign resultStage_mainTwoValidStream_payload = diffStage_mainTwoValidStream_s2mPipe_rData;
  assign diffStage_counterTwoValidStream_ready = (! diffStage_counterTwoValidStream_rValid);
  assign diffStage_counterTwoValidStream_s2mPipe_valid = (diffStage_counterTwoValidStream_valid || diffStage_counterTwoValidStream_rValid);
  assign diffStage_counterTwoValidStream_s2mPipe_payload = (diffStage_counterTwoValidStream_rValid ? diffStage_counterTwoValidStream_rData : diffStage_counterTwoValidStream_payload);
  always @(*) begin
    diffStage_counterTwoValidStream_s2mPipe_ready = resultStage_counterTwoValidStream_ready;
    if(when_Stream_l368_63) begin
      diffStage_counterTwoValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_63 = (! resultStage_counterTwoValidStream_valid);
  assign resultStage_counterTwoValidStream_valid = diffStage_counterTwoValidStream_s2mPipe_rValid;
  assign resultStage_counterTwoValidStream_payload = diffStage_counterTwoValidStream_s2mPipe_rData;
  assign diffStage_mainThreeValidStream_ready = (! diffStage_mainThreeValidStream_rValid);
  assign diffStage_mainThreeValidStream_s2mPipe_valid = (diffStage_mainThreeValidStream_valid || diffStage_mainThreeValidStream_rValid);
  assign diffStage_mainThreeValidStream_s2mPipe_payload = (diffStage_mainThreeValidStream_rValid ? diffStage_mainThreeValidStream_rData : diffStage_mainThreeValidStream_payload);
  always @(*) begin
    diffStage_mainThreeValidStream_s2mPipe_ready = resultStage_mainThreeValidStream_ready;
    if(when_Stream_l368_64) begin
      diffStage_mainThreeValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_64 = (! resultStage_mainThreeValidStream_valid);
  assign resultStage_mainThreeValidStream_valid = diffStage_mainThreeValidStream_s2mPipe_rValid;
  assign resultStage_mainThreeValidStream_payload = diffStage_mainThreeValidStream_s2mPipe_rData;
  assign diffStage_counterThreeValidStream_ready = (! diffStage_counterThreeValidStream_rValid);
  assign diffStage_counterThreeValidStream_s2mPipe_valid = (diffStage_counterThreeValidStream_valid || diffStage_counterThreeValidStream_rValid);
  assign diffStage_counterThreeValidStream_s2mPipe_payload = (diffStage_counterThreeValidStream_rValid ? diffStage_counterThreeValidStream_rData : diffStage_counterThreeValidStream_payload);
  always @(*) begin
    diffStage_counterThreeValidStream_s2mPipe_ready = resultStage_counterThreeValidStream_ready;
    if(when_Stream_l368_65) begin
      diffStage_counterThreeValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_65 = (! resultStage_counterThreeValidStream_valid);
  assign resultStage_counterThreeValidStream_valid = diffStage_counterThreeValidStream_s2mPipe_rValid;
  assign resultStage_counterThreeValidStream_payload = diffStage_counterThreeValidStream_s2mPipe_rData;
  assign diffStage_controlPipe_ready = diffStage_controlPipe_fork_io_input_ready;
  always @(*) begin
    CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin = diffStage_controlPipe_payload_isHorizontalMin;
    if(when_SuperResolutionPart3_l783) begin
      if(when_SuperResolutionPart3_l784) begin
        if(when_SuperResolutionPart3_l785) begin
          CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin = 1'b1;
        end else begin
          if(when_SuperResolutionPart3_l788) begin
            CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin = 1'b0;
          end else begin
            CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin = 1'b0;
          end
        end
      end else begin
        if(when_SuperResolutionPart3_l795) begin
          if(when_SuperResolutionPart3_l796) begin
            CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin = 1'b0;
          end else begin
            CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin = 1'b0;
          end
        end else begin
          if(when_SuperResolutionPart3_l803) begin
            if(when_SuperResolutionPart3_l804) begin
              CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin = 1'b1;
            end else begin
              CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin = 1'b0;
            end
          end else begin
            if(when_SuperResolutionPart3_l811) begin
              if(when_SuperResolutionPart3_l812) begin
                CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin = 1'b1;
              end else begin
                CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l819) begin
                CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin = 1'b0;
              end else begin
                if(when_SuperResolutionPart3_l822) begin
                  CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin = 1'b1;
                end else begin
                  if(when_SuperResolutionPart3_l825) begin
                    CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin = 1'b0;
                  end
                end
              end
            end
          end
        end
      end
    end
  end

  always @(*) begin
    CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff = diffStage_controlPipe_payload_minDiff;
    if(when_SuperResolutionPart3_l783) begin
      if(when_SuperResolutionPart3_l784) begin
        if(when_SuperResolutionPart3_l785) begin
          CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff = diffStage_controlPipe_payload_horizontalDiff;
        end else begin
          if(when_SuperResolutionPart3_l788) begin
            CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff = diffStage_controlPipe_payload_mainDiff;
          end else begin
            CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff = diffStage_controlPipe_payload_counterDiff;
          end
        end
      end else begin
        if(when_SuperResolutionPart3_l795) begin
          if(when_SuperResolutionPart3_l796) begin
            CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff = diffStage_controlPipe_payload_mainDiff;
          end else begin
            CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff = diffStage_controlPipe_payload_counterDiff;
          end
        end else begin
          if(when_SuperResolutionPart3_l803) begin
            if(when_SuperResolutionPart3_l804) begin
              CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff = diffStage_controlPipe_payload_horizontalDiff;
            end else begin
              CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff = diffStage_controlPipe_payload_counterDiff;
            end
          end else begin
            if(when_SuperResolutionPart3_l811) begin
              if(when_SuperResolutionPart3_l812) begin
                CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff = diffStage_controlPipe_payload_horizontalDiff;
              end else begin
                CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff = diffStage_controlPipe_payload_mainDiff;
              end
            end else begin
              if(when_SuperResolutionPart3_l819) begin
                CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff = diffStage_controlPipe_payload_counterDiff;
              end else begin
                if(when_SuperResolutionPart3_l822) begin
                  CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff = diffStage_controlPipe_payload_horizontalDiff;
                end else begin
                  if(when_SuperResolutionPart3_l825) begin
                    CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff = diffStage_controlPipe_payload_mainDiff;
                  end
                end
              end
            end
          end
        end
      end
    end
  end

  assign when_SuperResolutionPart3_l783 = (! diffStage_controlPipe_payload_finalResult);
  assign when_SuperResolutionPart3_l784 = ((diffStage_controlPipe_payload_horizontalDirectionValid && diffStage_controlPipe_payload_mainDirectionValid) && diffStage_controlPipe_payload_counterDirectionValid);
  assign when_SuperResolutionPart3_l785 = ((diffStage_controlPipe_payload_horizontalDiff <= diffStage_controlPipe_payload_mainDiff) && (diffStage_controlPipe_payload_horizontalDiff <= diffStage_controlPipe_payload_counterDiff));
  assign when_SuperResolutionPart3_l788 = ((diffStage_controlPipe_payload_mainDiff < diffStage_controlPipe_payload_horizontalDiff) && (diffStage_controlPipe_payload_mainDiff <= diffStage_controlPipe_payload_counterDiff));
  assign when_SuperResolutionPart3_l796 = (diffStage_controlPipe_payload_mainDiff <= diffStage_controlPipe_payload_counterDiff);
  assign when_SuperResolutionPart3_l804 = (diffStage_controlPipe_payload_horizontalDiff <= diffStage_controlPipe_payload_counterDiff);
  assign when_SuperResolutionPart3_l812 = (diffStage_controlPipe_payload_horizontalDiff <= diffStage_controlPipe_payload_mainDiff);
  assign when_SuperResolutionPart3_l795 = (((! diffStage_controlPipe_payload_horizontalDirectionValid) && diffStage_controlPipe_payload_mainDirectionValid) && diffStage_controlPipe_payload_counterDirectionValid);
  assign when_SuperResolutionPart3_l803 = ((diffStage_controlPipe_payload_horizontalDirectionValid && (! diffStage_controlPipe_payload_mainDirectionValid)) && diffStage_controlPipe_payload_counterDirectionValid);
  assign when_SuperResolutionPart3_l811 = ((diffStage_controlPipe_payload_horizontalDirectionValid && diffStage_controlPipe_payload_mainDirectionValid) && (! diffStage_controlPipe_payload_counterDirectionValid));
  assign when_SuperResolutionPart3_l819 = (((! diffStage_controlPipe_payload_horizontalDirectionValid) && (! diffStage_controlPipe_payload_mainDirectionValid)) && diffStage_controlPipe_payload_counterDirectionValid);
  assign when_SuperResolutionPart3_l822 = ((diffStage_controlPipe_payload_horizontalDirectionValid && (! diffStage_controlPipe_payload_mainDirectionValid)) && (! diffStage_controlPipe_payload_counterDirectionValid));
  assign when_SuperResolutionPart3_l825 = (((! diffStage_controlPipe_payload_horizontalDirectionValid) && diffStage_controlPipe_payload_mainDirectionValid) && (! diffStage_controlPipe_payload_counterDirectionValid));
  assign resultStage_controlPipeBeforePipe_valid = diffStage_controlPipe_fork_io_outputs_0_valid;
  assign resultStage_controlPipeBeforePipe_payload_frameStart = diffStage_controlPipe_payload_frameStart;
  assign resultStage_controlPipeBeforePipe_payload_rowEnd = diffStage_controlPipe_payload_rowEnd;
  assign resultStage_controlPipeBeforePipe_payload_pipeValid = diffStage_controlPipe_payload_pipeValid;
  assign resultStage_controlPipeBeforePipe_payload_firstRow = diffStage_controlPipe_payload_firstRow;
  assign resultStage_controlPipeBeforePipe_payload_lastRow = diffStage_controlPipe_payload_lastRow;
  assign resultStage_controlPipeBeforePipe_payload_finalResult = diffStage_controlPipe_payload_finalResult;
  assign resultStage_controlPipeBeforePipe_payload_mainCompare = diffStage_controlPipe_payload_mainCompare;
  assign resultStage_controlPipeBeforePipe_payload_counterCompare = diffStage_controlPipe_payload_counterCompare;
  assign resultStage_controlPipeBeforePipe_payload_horizontalCompare = diffStage_controlPipe_payload_horizontalCompare;
  assign resultStage_controlPipeBeforePipe_payload_verticalCompare = diffStage_controlPipe_payload_verticalCompare;
  assign resultStage_controlPipeBeforePipe_payload_mainDiff = diffStage_controlPipe_payload_mainDiff;
  assign resultStage_controlPipeBeforePipe_payload_counterDiff = diffStage_controlPipe_payload_counterDiff;
  assign resultStage_controlPipeBeforePipe_payload_horizontalDiff = diffStage_controlPipe_payload_horizontalDiff;
  assign resultStage_controlPipeBeforePipe_payload_verticalDiff = diffStage_controlPipe_payload_verticalDiff;
  assign resultStage_controlPipeBeforePipe_payload_isHorizontalMin = CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin;
  assign resultStage_controlPipeBeforePipe_payload_minDiff = CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff;
  assign resultStage_controlPipeBeforePipe_payload_currentPosition = diffStage_controlPipe_payload_currentPosition;
  assign resultStage_controlPipeBeforePipe_payload_nextPosition = diffStage_controlPipe_payload_nextPosition;
  assign resultStage_controlPipeBeforePipe_payload_horizontalDirectionValid = diffStage_controlPipe_payload_horizontalDirectionValid;
  assign resultStage_controlPipeBeforePipe_payload_verticalDirectionValid = diffStage_controlPipe_payload_verticalDirectionValid;
  assign resultStage_controlPipeBeforePipe_payload_mainDirectionValid = diffStage_controlPipe_payload_mainDirectionValid;
  assign resultStage_controlPipeBeforePipe_payload_counterDirectionValid = diffStage_controlPipe_payload_counterDirectionValid;
  assign resultStage_controlPipeBeforePipe_payload_inValidMinDiff = diffStage_controlPipe_payload_inValidMinDiff;
  assign resultStage_controlPipeBeforePipe_ready = (! resultStage_controlPipeBeforePipe_rValid);
  assign resultStage_controlPipeBeforePipe_s2mPipe_valid = (resultStage_controlPipeBeforePipe_valid || resultStage_controlPipeBeforePipe_rValid);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_frameStart = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_frameStart : resultStage_controlPipeBeforePipe_payload_frameStart);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_rowEnd = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_rowEnd : resultStage_controlPipeBeforePipe_payload_rowEnd);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_pipeValid = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_pipeValid : resultStage_controlPipeBeforePipe_payload_pipeValid);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_firstRow = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_firstRow : resultStage_controlPipeBeforePipe_payload_firstRow);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_lastRow = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_lastRow : resultStage_controlPipeBeforePipe_payload_lastRow);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_finalResult = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_finalResult : resultStage_controlPipeBeforePipe_payload_finalResult);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_mainCompare = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_mainCompare : resultStage_controlPipeBeforePipe_payload_mainCompare);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_counterCompare = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_counterCompare : resultStage_controlPipeBeforePipe_payload_counterCompare);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_horizontalCompare = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_horizontalCompare : resultStage_controlPipeBeforePipe_payload_horizontalCompare);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_verticalCompare = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_verticalCompare : resultStage_controlPipeBeforePipe_payload_verticalCompare);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_mainDiff = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_mainDiff : resultStage_controlPipeBeforePipe_payload_mainDiff);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_counterDiff = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_counterDiff : resultStage_controlPipeBeforePipe_payload_counterDiff);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_horizontalDiff = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_horizontalDiff : resultStage_controlPipeBeforePipe_payload_horizontalDiff);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_verticalDiff = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_verticalDiff : resultStage_controlPipeBeforePipe_payload_verticalDiff);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_isHorizontalMin = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_isHorizontalMin : resultStage_controlPipeBeforePipe_payload_isHorizontalMin);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_minDiff = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_minDiff : resultStage_controlPipeBeforePipe_payload_minDiff);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_currentPosition = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_currentPosition : resultStage_controlPipeBeforePipe_payload_currentPosition);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_nextPosition = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_nextPosition : resultStage_controlPipeBeforePipe_payload_nextPosition);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_horizontalDirectionValid = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_horizontalDirectionValid : resultStage_controlPipeBeforePipe_payload_horizontalDirectionValid);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_verticalDirectionValid = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_verticalDirectionValid : resultStage_controlPipeBeforePipe_payload_verticalDirectionValid);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_mainDirectionValid = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_mainDirectionValid : resultStage_controlPipeBeforePipe_payload_mainDirectionValid);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_counterDirectionValid = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_counterDirectionValid : resultStage_controlPipeBeforePipe_payload_counterDirectionValid);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_inValidMinDiff = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_inValidMinDiff : resultStage_controlPipeBeforePipe_payload_inValidMinDiff);
  always @(*) begin
    resultStage_controlPipeBeforePipe_s2mPipe_ready = resultStage_controlPipe_ready;
    if(when_Stream_l368_66) begin
      resultStage_controlPipeBeforePipe_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_66 = (! resultStage_controlPipe_valid);
  assign resultStage_controlPipe_valid = resultStage_controlPipeBeforePipe_s2mPipe_rValid;
  assign resultStage_controlPipe_payload_frameStart = resultStage_controlPipeBeforePipe_s2mPipe_rData_frameStart;
  assign resultStage_controlPipe_payload_rowEnd = resultStage_controlPipeBeforePipe_s2mPipe_rData_rowEnd;
  assign resultStage_controlPipe_payload_pipeValid = resultStage_controlPipeBeforePipe_s2mPipe_rData_pipeValid;
  assign resultStage_controlPipe_payload_firstRow = resultStage_controlPipeBeforePipe_s2mPipe_rData_firstRow;
  assign resultStage_controlPipe_payload_lastRow = resultStage_controlPipeBeforePipe_s2mPipe_rData_lastRow;
  assign resultStage_controlPipe_payload_finalResult = resultStage_controlPipeBeforePipe_s2mPipe_rData_finalResult;
  assign resultStage_controlPipe_payload_mainCompare = resultStage_controlPipeBeforePipe_s2mPipe_rData_mainCompare;
  assign resultStage_controlPipe_payload_counterCompare = resultStage_controlPipeBeforePipe_s2mPipe_rData_counterCompare;
  assign resultStage_controlPipe_payload_horizontalCompare = resultStage_controlPipeBeforePipe_s2mPipe_rData_horizontalCompare;
  assign resultStage_controlPipe_payload_verticalCompare = resultStage_controlPipeBeforePipe_s2mPipe_rData_verticalCompare;
  assign resultStage_controlPipe_payload_mainDiff = resultStage_controlPipeBeforePipe_s2mPipe_rData_mainDiff;
  assign resultStage_controlPipe_payload_counterDiff = resultStage_controlPipeBeforePipe_s2mPipe_rData_counterDiff;
  assign resultStage_controlPipe_payload_horizontalDiff = resultStage_controlPipeBeforePipe_s2mPipe_rData_horizontalDiff;
  assign resultStage_controlPipe_payload_verticalDiff = resultStage_controlPipeBeforePipe_s2mPipe_rData_verticalDiff;
  assign resultStage_controlPipe_payload_isHorizontalMin = resultStage_controlPipeBeforePipe_s2mPipe_rData_isHorizontalMin;
  assign resultStage_controlPipe_payload_minDiff = resultStage_controlPipeBeforePipe_s2mPipe_rData_minDiff;
  assign resultStage_controlPipe_payload_currentPosition = resultStage_controlPipeBeforePipe_s2mPipe_rData_currentPosition;
  assign resultStage_controlPipe_payload_nextPosition = resultStage_controlPipeBeforePipe_s2mPipe_rData_nextPosition;
  assign resultStage_controlPipe_payload_horizontalDirectionValid = resultStage_controlPipeBeforePipe_s2mPipe_rData_horizontalDirectionValid;
  assign resultStage_controlPipe_payload_verticalDirectionValid = resultStage_controlPipeBeforePipe_s2mPipe_rData_verticalDirectionValid;
  assign resultStage_controlPipe_payload_mainDirectionValid = resultStage_controlPipeBeforePipe_s2mPipe_rData_mainDirectionValid;
  assign resultStage_controlPipe_payload_counterDirectionValid = resultStage_controlPipeBeforePipe_s2mPipe_rData_counterDirectionValid;
  assign resultStage_controlPipe_payload_inValidMinDiff = resultStage_controlPipeBeforePipe_s2mPipe_rData_inValidMinDiff;
  assign resultStage_pixelStream_valid = diffStage_controlPipe_fork_io_outputs_1_valid;
  always @(*) begin
    resultStage_pixelStream_payload = 8'h0;
    if(diffStage_controlPipe_payload_finalResult) begin
      if(when_SuperResolutionPart3_l840) begin
        resultStage_pixelStream_payload = diffStage_mainOnePixelStream_payload;
      end else begin
        if(when_SuperResolutionPart3_l841) begin
          resultStage_pixelStream_payload = diffStage_mainTwoPixelStream_payload;
        end else begin
          if(when_SuperResolutionPart3_l842) begin
            resultStage_pixelStream_payload = diffStage_mainThreePixelStream_payload;
          end else begin
            if(diffStage_controlPipe_payload_verticalDirectionValid) begin
              if(inValidMinDiff) begin
                if(when_SuperResolutionPart3_l846) begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload[7:0];
                end else begin
                  if(when_SuperResolutionPart3_l847) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_2[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_4[7:0];
                  end
                end
              end else begin
                if(when_SuperResolutionPart3_l850) begin
                  resultStage_pixelStream_payload = candidatePixel;
                end else begin
                  if(when_SuperResolutionPart3_l851) begin
                    if(isHorizontalDirection) begin
                      resultStage_pixelStream_payload = candidatePixel;
                    end else begin
                      if(when_SuperResolutionPart3_l854) begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_6[7:0];
                      end else begin
                        if(when_SuperResolutionPart3_l855) begin
                          resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_8[7:0];
                        end else begin
                          resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_10[7:0];
                        end
                      end
                    end
                  end else begin
                    if(when_SuperResolutionPart3_l860) begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_12[7:0];
                    end else begin
                      if(when_SuperResolutionPart3_l861) begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_14[7:0];
                      end else begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_16[7:0];
                      end
                    end
                  end
                end
              end
            end else begin
              resultStage_pixelStream_payload = candidatePixel;
            end
          end
        end
      end
    end else begin
      if(when_SuperResolutionPart3_l869) begin
        if(when_SuperResolutionPart3_l870) begin
          if(when_SuperResolutionPart3_l871) begin
            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_18[7:0];
          end else begin
            if(when_SuperResolutionPart3_l872) begin
              resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_20[7:0];
            end else begin
              resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_22[7:0];
            end
          end
        end else begin
          if(when_SuperResolutionPart3_l874) begin
            if(when_SuperResolutionPart3_l875) begin
              if(when_SuperResolutionPart3_l876) begin
                if(diffStage_controlPipe_payload_firstRow) begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_24[7:0];
                end else begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_26[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_28[7:0];
                  end
                end
              end else begin
                if(diffStage_controlPipe_payload_lastRow) begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_30[7:0];
                end else begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_32[7:0];
                end
              end
            end else begin
              if(when_SuperResolutionPart3_l884) begin
                if(when_SuperResolutionPart3_l885) begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_34[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_36[7:0];
                  end
                end else begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_38[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_40[7:0];
                  end
                end
              end else begin
                if(when_SuperResolutionPart3_l893) begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_42[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_44[7:0];
                  end
                end else begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_46[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_48[7:0];
                  end
                end
              end
            end
          end else begin
            if(when_SuperResolutionPart3_l902) begin
              if(when_SuperResolutionPart3_l903) begin
                if(diffStage_controlPipe_payload_firstRow) begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_50[7:0];
                end else begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_52[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_54[7:0];
                  end
                end
              end else begin
                if(diffStage_controlPipe_payload_lastRow) begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_56[7:0];
                end else begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_58[7:0];
                end
              end
            end else begin
              if(when_SuperResolutionPart3_l911) begin
                if(when_SuperResolutionPart3_l912) begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_60[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_62[7:0];
                  end
                end else begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_64[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_66[7:0];
                  end
                end
              end else begin
                if(when_SuperResolutionPart3_l920) begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_68[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_70[7:0];
                  end
                end else begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_72[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_74[7:0];
                  end
                end
              end
            end
          end
        end
      end else begin
        if(when_SuperResolutionPart3_l929) begin
          if(when_SuperResolutionPart3_l930) begin
            if(when_SuperResolutionPart3_l931) begin
              if(when_SuperResolutionPart3_l932) begin
                if(diffStage_controlPipe_payload_firstRow) begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_76[7:0];
                end else begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_78[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_80[7:0];
                  end
                end
              end else begin
                if(diffStage_controlPipe_payload_lastRow) begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_82[7:0];
                end else begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_84[7:0];
                end
              end
            end else begin
              if(when_SuperResolutionPart3_l940) begin
                if(when_SuperResolutionPart3_l941) begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_86[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_88[7:0];
                  end
                end else begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_90[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_92[7:0];
                  end
                end
              end else begin
                if(when_SuperResolutionPart3_l949) begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_94[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_96[7:0];
                  end
                end else begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_98[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_100[7:0];
                  end
                end
              end
            end
          end else begin
            if(when_SuperResolutionPart3_l958) begin
              if(when_SuperResolutionPart3_l959) begin
                if(diffStage_controlPipe_payload_firstRow) begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_102[7:0];
                end else begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_104[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_106[7:0];
                  end
                end
              end else begin
                if(diffStage_controlPipe_payload_lastRow) begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_108[7:0];
                end else begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_110[7:0];
                end
              end
            end else begin
              if(when_SuperResolutionPart3_l967) begin
                if(when_SuperResolutionPart3_l968) begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_112[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_114[7:0];
                  end
                end else begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_116[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_118[7:0];
                  end
                end
              end else begin
                if(when_SuperResolutionPart3_l976) begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_120[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_122[7:0];
                  end
                end else begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_124[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_126[7:0];
                  end
                end
              end
            end
          end
        end else begin
          if(when_SuperResolutionPart3_l985) begin
            if(when_SuperResolutionPart3_l986) begin
              if(when_SuperResolutionPart3_l987) begin
                resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_128[7:0];
              end else begin
                if(when_SuperResolutionPart3_l988) begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_130[7:0];
                end else begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_132[7:0];
                end
              end
            end else begin
              if(when_SuperResolutionPart3_l991) begin
                if(when_SuperResolutionPart3_l992) begin
                  if(diffStage_controlPipe_payload_firstRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_134[7:0];
                  end else begin
                    if(diffStage_controlPipe_payload_lastRow) begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_136[7:0];
                    end else begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_138[7:0];
                    end
                  end
                end else begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_140[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_142[7:0];
                  end
                end
              end else begin
                if(when_SuperResolutionPart3_l1000) begin
                  if(when_SuperResolutionPart3_l1001) begin
                    if(diffStage_controlPipe_payload_lastRow) begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_144[7:0];
                    end else begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_146[7:0];
                    end
                  end else begin
                    if(diffStage_controlPipe_payload_lastRow) begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_148[7:0];
                    end else begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_150[7:0];
                    end
                  end
                end else begin
                  if(when_SuperResolutionPart3_l1009) begin
                    if(diffStage_controlPipe_payload_lastRow) begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_152[7:0];
                    end else begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_154[7:0];
                    end
                  end else begin
                    if(diffStage_controlPipe_payload_lastRow) begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_156[7:0];
                    end else begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_158[7:0];
                    end
                  end
                end
              end
            end
          end else begin
            if(when_SuperResolutionPart3_l1018) begin
              if(when_SuperResolutionPart3_l1019) begin
                if(when_SuperResolutionPart3_l1020) begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_160[7:0];
                end else begin
                  if(when_SuperResolutionPart3_l1021) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_162[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_164[7:0];
                  end
                end
              end else begin
                if(when_SuperResolutionPart3_l1024) begin
                  if(when_SuperResolutionPart3_l1025) begin
                    if(diffStage_controlPipe_payload_firstRow) begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_166[7:0];
                    end else begin
                      if(diffStage_controlPipe_payload_lastRow) begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_168[7:0];
                      end else begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_170[7:0];
                      end
                    end
                  end else begin
                    if(diffStage_controlPipe_payload_lastRow) begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_172[7:0];
                    end else begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_174[7:0];
                    end
                  end
                end else begin
                  if(when_SuperResolutionPart3_l1033) begin
                    if(when_SuperResolutionPart3_l1034) begin
                      if(diffStage_controlPipe_payload_lastRow) begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_176[7:0];
                      end else begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_178[7:0];
                      end
                    end else begin
                      if(diffStage_controlPipe_payload_lastRow) begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_180[7:0];
                      end else begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_182[7:0];
                      end
                    end
                  end else begin
                    if(when_SuperResolutionPart3_l1042) begin
                      if(diffStage_controlPipe_payload_lastRow) begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_184[7:0];
                      end else begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_186[7:0];
                      end
                    end else begin
                      if(diffStage_controlPipe_payload_lastRow) begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_188[7:0];
                      end else begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_190[7:0];
                      end
                    end
                  end
                end
              end
            end else begin
              if(when_SuperResolutionPart3_l1051) begin
                if(when_SuperResolutionPart3_l1052) begin
                  if(when_SuperResolutionPart3_l1053) begin
                    if(diffStage_controlPipe_payload_firstRow) begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_192[7:0];
                    end else begin
                      if(diffStage_controlPipe_payload_lastRow) begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_194[7:0];
                      end else begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_196[7:0];
                      end
                    end
                  end else begin
                    if(diffStage_controlPipe_payload_lastRow) begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_198[7:0];
                    end else begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_200[7:0];
                    end
                  end
                end else begin
                  if(when_SuperResolutionPart3_l1061) begin
                    if(when_SuperResolutionPart3_l1062) begin
                      if(diffStage_controlPipe_payload_lastRow) begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_202[7:0];
                      end else begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_204[7:0];
                      end
                    end else begin
                      if(diffStage_controlPipe_payload_lastRow) begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_206[7:0];
                      end else begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_208[7:0];
                      end
                    end
                  end else begin
                    if(when_SuperResolutionPart3_l1070) begin
                      if(diffStage_controlPipe_payload_lastRow) begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_210[7:0];
                      end else begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_212[7:0];
                      end
                    end else begin
                      if(diffStage_controlPipe_payload_lastRow) begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_214[7:0];
                      end else begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_216[7:0];
                      end
                    end
                  end
                end
              end else begin
                if(when_SuperResolutionPart3_l1078) begin
                  if(when_SuperResolutionPart3_l1079) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_218[7:0];
                  end else begin
                    if(when_SuperResolutionPart3_l1080) begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_220[7:0];
                    end else begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_222[7:0];
                    end
                  end
                end else begin
                  if(when_SuperResolutionPart3_l1082) begin
                    if(when_SuperResolutionPart3_l1083) begin
                      if(when_SuperResolutionPart3_l1084) begin
                        if(diffStage_controlPipe_payload_firstRow) begin
                          resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_224[7:0];
                        end else begin
                          if(diffStage_controlPipe_payload_lastRow) begin
                            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_226[7:0];
                          end else begin
                            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_228[7:0];
                          end
                        end
                      end else begin
                        if(diffStage_controlPipe_payload_lastRow) begin
                          resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_230[7:0];
                        end else begin
                          resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_232[7:0];
                        end
                      end
                    end else begin
                      if(when_SuperResolutionPart3_l1092) begin
                        if(when_SuperResolutionPart3_l1093) begin
                          if(diffStage_controlPipe_payload_lastRow) begin
                            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_234[7:0];
                          end else begin
                            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_236[7:0];
                          end
                        end else begin
                          if(diffStage_controlPipe_payload_lastRow) begin
                            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_238[7:0];
                          end else begin
                            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_240[7:0];
                          end
                        end
                      end else begin
                        if(when_SuperResolutionPart3_l1101) begin
                          if(diffStage_controlPipe_payload_lastRow) begin
                            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_242[7:0];
                          end else begin
                            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_244[7:0];
                          end
                        end else begin
                          if(diffStage_controlPipe_payload_lastRow) begin
                            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_246[7:0];
                          end else begin
                            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_248[7:0];
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
  end

  assign when_SuperResolutionPart3_l840 = ((diffStage_controlPipe_payload_currentPosition == 2'b00) && diffStage_mainOneValidStream_payload);
  assign when_SuperResolutionPart3_l846 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l847 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l850 = (minDiff < diffStage_controlPipe_payload_verticalDiff);
  assign when_SuperResolutionPart3_l854 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l855 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l860 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l861 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l851 = (diffStage_controlPipe_payload_verticalDiff == minDiff);
  assign when_SuperResolutionPart3_l841 = ((diffStage_controlPipe_payload_currentPosition == 2'b01) && diffStage_mainTwoValidStream_payload);
  assign when_SuperResolutionPart3_l842 = ((diffStage_controlPipe_payload_currentPosition == 2'b10) && diffStage_mainThreeValidStream_payload);
  assign when_SuperResolutionPart3_l869 = ((diffStage_controlPipe_payload_horizontalDirectionValid && diffStage_controlPipe_payload_mainDirectionValid) && diffStage_controlPipe_payload_counterDirectionValid);
  assign when_SuperResolutionPart3_l870 = ((diffStage_controlPipe_payload_horizontalDiff <= diffStage_controlPipe_payload_mainDiff) && (diffStage_controlPipe_payload_horizontalDiff <= diffStage_controlPipe_payload_counterDiff));
  assign when_SuperResolutionPart3_l871 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l872 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l875 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l876 = (diffStage_controlPipe_payload_nextPosition == 2'b01);
  assign when_SuperResolutionPart3_l885 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l893 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l884 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l902 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l903 = (diffStage_controlPipe_payload_nextPosition == 2'b01);
  assign when_SuperResolutionPart3_l912 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l920 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l911 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l874 = ((diffStage_controlPipe_payload_mainDiff < diffStage_controlPipe_payload_horizontalDiff) && (diffStage_controlPipe_payload_mainDiff <= diffStage_controlPipe_payload_counterDiff));
  assign when_SuperResolutionPart3_l930 = (diffStage_controlPipe_payload_mainDiff <= diffStage_controlPipe_payload_counterDiff);
  assign when_SuperResolutionPart3_l931 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l932 = (diffStage_controlPipe_payload_nextPosition == 2'b01);
  assign when_SuperResolutionPart3_l941 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l949 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l940 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l958 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l959 = (diffStage_controlPipe_payload_nextPosition == 2'b01);
  assign when_SuperResolutionPart3_l968 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l976 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l967 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l986 = (diffStage_controlPipe_payload_horizontalDiff <= diffStage_controlPipe_payload_counterDiff);
  assign when_SuperResolutionPart3_l987 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l988 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l991 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l992 = (diffStage_controlPipe_payload_nextPosition == 2'b01);
  assign when_SuperResolutionPart3_l1001 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l1009 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l1000 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l1019 = (diffStage_controlPipe_payload_horizontalDiff <= diffStage_controlPipe_payload_mainDiff);
  assign when_SuperResolutionPart3_l1020 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l1021 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l1024 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l1025 = (diffStage_controlPipe_payload_nextPosition == 2'b01);
  assign when_SuperResolutionPart3_l1034 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l1042 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l1033 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l1052 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l1053 = (diffStage_controlPipe_payload_nextPosition == 2'b01);
  assign when_SuperResolutionPart3_l1062 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l1070 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l1061 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l1079 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l1080 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l1083 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l1084 = (diffStage_controlPipe_payload_nextPosition == 2'b01);
  assign when_SuperResolutionPart3_l1093 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l1101 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l1092 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l929 = (((! diffStage_controlPipe_payload_horizontalDirectionValid) && diffStage_controlPipe_payload_mainDirectionValid) && diffStage_controlPipe_payload_counterDirectionValid);
  assign when_SuperResolutionPart3_l985 = ((diffStage_controlPipe_payload_horizontalDirectionValid && (! diffStage_controlPipe_payload_mainDirectionValid)) && diffStage_controlPipe_payload_counterDirectionValid);
  assign when_SuperResolutionPart3_l1018 = ((diffStage_controlPipe_payload_horizontalDirectionValid && diffStage_controlPipe_payload_mainDirectionValid) && (! diffStage_controlPipe_payload_counterDirectionValid));
  assign when_SuperResolutionPart3_l1051 = (((! diffStage_controlPipe_payload_horizontalDirectionValid) && (! diffStage_controlPipe_payload_mainDirectionValid)) && diffStage_controlPipe_payload_counterDirectionValid);
  assign when_SuperResolutionPart3_l1078 = ((diffStage_controlPipe_payload_horizontalDirectionValid && (! diffStage_controlPipe_payload_mainDirectionValid)) && (! diffStage_controlPipe_payload_counterDirectionValid));
  assign when_SuperResolutionPart3_l1082 = (((! diffStage_controlPipe_payload_horizontalDirectionValid) && diffStage_controlPipe_payload_mainDirectionValid) && (! diffStage_controlPipe_payload_counterDirectionValid));
  assign resultStage_pixelStream_ready = (! resultStage_pixelStream_rValid);
  assign resultStage_pixelStream_s2mPipe_valid = (resultStage_pixelStream_valid || resultStage_pixelStream_rValid);
  assign resultStage_pixelStream_s2mPipe_payload = (resultStage_pixelStream_rValid ? resultStage_pixelStream_rData : resultStage_pixelStream_payload);
  always @(*) begin
    resultStage_pixelStream_s2mPipe_ready = resultStage_resultStream_ready;
    if(when_Stream_l368_67) begin
      resultStage_pixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_67 = (! resultStage_resultStream_valid);
  assign resultStage_resultStream_valid = resultStage_pixelStream_s2mPipe_rValid;
  assign resultStage_resultStream_payload = resultStage_pixelStream_s2mPipe_rData;
  assign when_SuperResolutionPart3_l1115 = (! resultStage_controlPipeBeforePipe_payload_finalResult);
  assign diffStage_controlPipe_fire = (diffStage_controlPipe_valid && diffStage_controlPipe_ready);
  assign CICC1851_resultStage_mainOnePixelStream_ready_2 = (CICC1851_resultStage_mainOnePixelStream_ready && CICC1851_resultStage_mainOnePixelStream_ready_1);
  assign CICC1851_resultStage_mainOnePixelStream_ready = (((((((((((((resultStage_resultStream_valid && resultStage_mainOnePixelStream_valid) && resultStage_counterOnePixelStream_valid) && resultStage_mainTwoPixelStream_valid) && resultStage_counterTwoPixelStream_valid) && resultStage_mainThreePixelStream_valid) && resultStage_counterThreePixelStream_valid) && resultStage_mainOneValidStream_valid) && resultStage_counterOneValidStream_valid) && resultStage_mainTwoValidStream_valid) && resultStage_counterTwoValidStream_valid) && resultStage_mainThreeValidStream_valid) && resultStage_counterThreeValidStream_valid) && resultStage_controlPipe_valid);
  assign resultStage_resultStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_mainOnePixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_counterOnePixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_mainTwoPixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_counterTwoPixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_mainThreePixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_counterThreePixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_mainOneValidStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_counterOneValidStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_mainTwoValidStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_counterTwoValidStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_mainThreeValidStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_counterThreeValidStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_controlPipe_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign when_Stream_l438 = ((! resultStage_controlPipe_payload_pipeValid) || (! resultStage_controlPipe_payload_finalResult));
  always @(*) begin
    resultsJoin_valid = CICC1851_resultStage_mainOnePixelStream_ready;
    if(when_Stream_l438) begin
      resultsJoin_valid = 1'b0;
    end
  end

  always @(*) begin
    CICC1851_resultStage_mainOnePixelStream_ready_1 = resultsJoin_ready;
    if(when_Stream_l438) begin
      CICC1851_resultStage_mainOnePixelStream_ready_1 = 1'b1;
    end
  end

  assign pixelsStream_valid = resultsJoin_valid;
  assign resultsJoin_ready = pixelsStream_ready;
  assign pixelsStream_payload_pixel = resultStage_resultStream_payload;
  assign pixelsStream_payload_frameStart = resultStage_controlPipe_payload_frameStart;
  assign pixelsStream_payload_rowEnd = resultStage_controlPipe_payload_rowEnd;
  assign pixelsStream_ready = (! pixelsStream_rValid);
  assign pixelsStream_s2mPipe_valid = (pixelsStream_valid || pixelsStream_rValid);
  assign pixelsStream_s2mPipe_payload_pixel = (pixelsStream_rValid ? pixelsStream_rData_pixel : pixelsStream_payload_pixel);
  assign pixelsStream_s2mPipe_payload_frameStart = (pixelsStream_rValid ? pixelsStream_rData_frameStart : pixelsStream_payload_frameStart);
  assign pixelsStream_s2mPipe_payload_rowEnd = (pixelsStream_rValid ? pixelsStream_rData_rowEnd : pixelsStream_payload_rowEnd);
  always @(*) begin
    pixelsStream_s2mPipe_ready = pixelsStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_68) begin
      pixelsStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_68 = (! pixelsStream_s2mPipe_m2sPipe_valid);
  assign pixelsStream_s2mPipe_m2sPipe_valid = pixelsStream_s2mPipe_rValid;
  assign pixelsStream_s2mPipe_m2sPipe_payload_pixel = pixelsStream_s2mPipe_rData_pixel;
  assign pixelsStream_s2mPipe_m2sPipe_payload_frameStart = pixelsStream_s2mPipe_rData_frameStart;
  assign pixelsStream_s2mPipe_m2sPipe_payload_rowEnd = pixelsStream_s2mPipe_rData_rowEnd;
  assign pixelsStream_s2mPipe_m2sPipe_ready = pixelsOut_ready;
  assign controlStateMachine_wantExit = 1'b0;
  always @(*) begin
    controlStateMachine_wantStart = 1'b0;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_5_HOLD : begin
      end
      controlStateMachine_enumDef_5_PASS : begin
      end
      controlStateMachine_enumDef_5_EXTRA : begin
      end
      default : begin
        controlStateMachine_wantStart = 1'b1;
      end
    endcase
  end

  assign controlStateMachine_wantKill = 1'b0;
  always @(*) begin
    controlStateMachine_stateNext = controlStateMachine_stateReg;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_5_HOLD : begin
        if(passPixels_fire_13) begin
          if(when_SuperResolutionPart3_l1158) begin
            controlStateMachine_stateNext = controlStateMachine_enumDef_5_PASS;
          end
        end
      end
      controlStateMachine_enumDef_5_PASS : begin
        if(controlStream_fire) begin
          controlStateMachine_stateNext = controlStateMachine_enumDef_5_EXTRA;
        end
      end
      controlStateMachine_enumDef_5_EXTRA : begin
        if(controlStream_fire_1) begin
          if(writeDone) begin
            if(when_SuperResolutionPart3_l1199) begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_5_HOLD;
            end else begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_5_PASS;
            end
          end else begin
            if(outReachRowEnd) begin
              if(when_SuperResolutionPart3_l1202) begin
                controlStateMachine_stateNext = controlStateMachine_enumDef_5_PASS;
              end else begin
                controlStateMachine_stateNext = controlStateMachine_enumDef_5_HOLD;
              end
            end else begin
              if(when_SuperResolutionPart3_l1205) begin
                controlStateMachine_stateNext = controlStateMachine_enumDef_5_PASS;
              end else begin
                controlStateMachine_stateNext = controlStateMachine_enumDef_5_HOLD;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
    if(controlStateMachine_wantStart) begin
      controlStateMachine_stateNext = controlStateMachine_enumDef_5_HOLD;
    end
    if(controlStateMachine_wantKill) begin
      controlStateMachine_stateNext = controlStateMachine_enumDef_5_BOOT;
    end
  end

  assign passPixels_fire_13 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart3_l1158 = ((outRowCount_value < bufferRowCount_value) && (outPixelAddr_value < bufferWAddr_value));
  assign controlStream_fire = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart3_l1168 = (outPixelAddr_value == 12'h0);
  assign when_SuperResolutionPart3_l1188 = (outRowCount_value == 12'h0);
  assign controlStream_fire_1 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart3_l1199 = (outReachFinalRow && outReachRowEnd);
  assign passPixels_fire_14 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart3_l1202 = (((bufferRowCount_value == CICC1851_when_SuperResolutionPart3_l1202) || (12'h001 < bufferWAddr_value)) || ((bufferWAddr_value == 12'h001) && passPixels_fire_14));
  assign passPixels_fire_15 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart3_l1205 = (((CICC1851_when_SuperResolutionPart3_l1205 < bufferRowCount_value) || ((bufferWAddr_value == CICC1851_when_SuperResolutionPart3_l1205_1) && passPixels_fire_15)) || (CICC1851_when_SuperResolutionPart3_l1205_2 < bufferWAddr_value));
  assign when_SuperResolutionPart3_l1217 = (outRowCount_value == 12'h0);
  assign controlStream_fire_2 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart3_l1220 = (frameStart && controlStream_fire_2);
  assign controlStream_fire_3 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart3_l1223 = (controlStream_fire_3 && (CICC1851_when_SuperResolutionPart3_l1223 == CICC1851_when_SuperResolutionPart3_l1223_1));
  assign controlStream_fire_4 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart3_l1224 = ((outReachRowEnd && (CICC1851_when_SuperResolutionPart3_l1224 == CICC1851_when_SuperResolutionPart3_l1224_1)) && controlStream_fire_4);
  assign controlStream_fire_5 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart3_l1226 = (controlStream_fire_5 && outReachRowEnd);
  assign controlStream_fire_6 = (controlStream_valid && controlStream_ready);
  assign controlStream_fire_7 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart3_l1247 = (controlStream_payload_rowEnd && controlStream_fire_7);
  assign when_SuperResolutionPart3_l1248 = (outRowCount_value != 12'h0);
  assign when_SuperResolutionPart3_l1250 = (currentRowBuffer == 2'b10);
  assign when_SuperResolutionPart3_l1252 = (nextRowBuffer == 2'b10);
  always @(posedge clk or negedge resetn) begin
    if(!resetn) begin
      inpThreeDone <= 1'b0;
      readDone <= 1'b0;
      startRead <= 1'b0;
      frameStart <= 1'b0;
      inpThreshold <= 8'h80;
      bmpWidth <= 10'h3c0;
      bmpHeight <= 10'h21c;
      holdBuffer <= 1'b0;
      writeDone <= 1'b0;
      bufferRowCount_value <= 12'h0;
      bufferEnable <= 1'b0;
      bufferSwitch <= 2'b00;
      nextRowBuffer <= 2'b01;
      currentRowBuffer <= 2'b00;
      bufferReuse <= 1'b0;
      bufferWAddr_value <= 12'h0;
      outPixelAddr_value <= 12'h0;
      outRowCount_value <= 12'h0;
      alreadySendRow_value <= 12'h0;
      alreadySendCountInRow_value <= 12'h0;
      alreadyReachRowEnd <= 1'b0;
      alreadyReachFinalRow <= 1'b0;
      outReachRowEnd <= 1'b0;
      outReachFinalRow <= 1'b0;
      bufferReachRowEnd <= 1'b0;
      bufferReachFinalRow <= 1'b0;
      minDiff <= 8'h0;
      candidatePixel <= 8'h0;
      isHorizontalDirection <= 1'b0;
      inValidMinDiff <= 1'b0;
      pixelsIn_rValid <= 1'b0;
      pixelsIn_s2mPipe_rValid <= 1'b0;
      mainPixelAddrOneStream_rValid <= 1'b0;
      mainPixelAddrOneStream_s2mPipe_rValid <= 1'b0;
      CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_mainOnePixelStream_valid <= 1'b0;
      counterPixelAddrOneStream_rValid <= 1'b0;
      counterPixelAddrOneStream_s2mPipe_rValid <= 1'b0;
      CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_counterOnePixelStream_valid <= 1'b0;
      mainPixelAddrTwoStream_rValid <= 1'b0;
      mainPixelAddrTwoStream_s2mPipe_rValid <= 1'b0;
      CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_mainTwoPixelStream_valid <= 1'b0;
      counterPixelAddrTwoStream_rValid <= 1'b0;
      counterPixelAddrTwoStream_s2mPipe_rValid <= 1'b0;
      CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_counterTwoPixelStream_valid <= 1'b0;
      mainPixelAddrThreeStream_rValid <= 1'b0;
      mainPixelAddrThreeStream_s2mPipe_rValid <= 1'b0;
      CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_mainThreePixelStream_valid <= 1'b0;
      counterPixelAddrThreeStream_rValid <= 1'b0;
      counterPixelAddrThreeStream_s2mPipe_rValid <= 1'b0;
      CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_counterThreePixelStream_valid <= 1'b0;
      mainValidAddrOneStream_rValid <= 1'b0;
      mainValidAddrOneStream_s2mPipe_rValid <= 1'b0;
      CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_mainOneValidStream_valid <= 1'b0;
      counterValidAddrOneStream_rValid <= 1'b0;
      counterValidAddrOneStream_s2mPipe_rValid <= 1'b0;
      CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_counterOneValidStream_valid <= 1'b0;
      mainValidAddrTwoStream_rValid <= 1'b0;
      mainValidAddrTwoStream_s2mPipe_rValid <= 1'b0;
      CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_mainTwoValidStream_valid <= 1'b0;
      counterValidAddrTwoStream_rValid <= 1'b0;
      counterValidAddrTwoStream_s2mPipe_rValid <= 1'b0;
      CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_counterTwoValidStream_valid <= 1'b0;
      mainValidAddrThreeStream_rValid <= 1'b0;
      mainValidAddrThreeStream_s2mPipe_rValid <= 1'b0;
      CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_mainThreeValidStream_valid <= 1'b0;
      counterValidAddrThreeStream_rValid <= 1'b0;
      counterValidAddrThreeStream_s2mPipe_rValid <= 1'b0;
      CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_counterThreeValidStream_valid <= 1'b0;
      controlStream_rValid <= 1'b0;
      controlStream_s2mPipe_rValid <= 1'b0;
      controlStream_s2mPipe_m2sPipe_rValid <= 1'b0;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rValid <= 1'b0;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rValid <= 1'b0;
      readStage_mainOnePixelStream_rValid <= 1'b0;
      readStage_mainOnePixelStream_s2mPipe_rValid <= 1'b0;
      readStage_counterOnePixelStream_rValid <= 1'b0;
      readStage_counterOnePixelStream_s2mPipe_rValid <= 1'b0;
      readStage_mainTwoPixelStream_rValid <= 1'b0;
      readStage_mainTwoPixelStream_s2mPipe_rValid <= 1'b0;
      readStage_counterTwoPixelStream_rValid <= 1'b0;
      readStage_counterTwoPixelStream_s2mPipe_rValid <= 1'b0;
      readStage_mainThreePixelStream_rValid <= 1'b0;
      readStage_mainThreePixelStream_s2mPipe_rValid <= 1'b0;
      readStage_counterThreePixelStream_rValid <= 1'b0;
      readStage_counterThreePixelStream_s2mPipe_rValid <= 1'b0;
      readStage_mainOneValidStream_rValid <= 1'b0;
      readStage_mainOneValidStream_s2mPipe_rValid <= 1'b0;
      readStage_counterOneValidStream_rValid <= 1'b0;
      readStage_counterOneValidStream_s2mPipe_rValid <= 1'b0;
      readStage_mainTwoValidStream_rValid <= 1'b0;
      readStage_mainTwoValidStream_s2mPipe_rValid <= 1'b0;
      readStage_counterTwoValidStream_rValid <= 1'b0;
      readStage_counterTwoValidStream_s2mPipe_rValid <= 1'b0;
      readStage_mainThreeValidStream_rValid <= 1'b0;
      readStage_mainThreeValidStream_s2mPipe_rValid <= 1'b0;
      readStage_counterThreeValidStream_rValid <= 1'b0;
      readStage_counterThreeValidStream_s2mPipe_rValid <= 1'b0;
      readStage_controlPipe_translated_rValid <= 1'b0;
      readStage_controlPipe_translated_s2mPipe_rValid <= 1'b0;
      compareStage_mainOnePixelStream_rValid <= 1'b0;
      compareStage_mainOnePixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_counterOnePixelStream_rValid <= 1'b0;
      compareStage_counterOnePixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_mainTwoPixelStream_rValid <= 1'b0;
      compareStage_mainTwoPixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_counterTwoPixelStream_rValid <= 1'b0;
      compareStage_counterTwoPixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_mainThreePixelStream_rValid <= 1'b0;
      compareStage_mainThreePixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_counterThreePixelStream_rValid <= 1'b0;
      compareStage_counterThreePixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_mainOneValidStream_rValid <= 1'b0;
      compareStage_mainOneValidStream_s2mPipe_rValid <= 1'b0;
      compareStage_counterOneValidStream_rValid <= 1'b0;
      compareStage_counterOneValidStream_s2mPipe_rValid <= 1'b0;
      compareStage_mainTwoValidStream_rValid <= 1'b0;
      compareStage_mainTwoValidStream_s2mPipe_rValid <= 1'b0;
      compareStage_counterTwoValidStream_rValid <= 1'b0;
      compareStage_counterTwoValidStream_s2mPipe_rValid <= 1'b0;
      compareStage_mainThreeValidStream_rValid <= 1'b0;
      compareStage_mainThreeValidStream_s2mPipe_rValid <= 1'b0;
      compareStage_counterThreeValidStream_rValid <= 1'b0;
      compareStage_counterThreeValidStream_s2mPipe_rValid <= 1'b0;
      compareStage_controlPipe_translated_rValid <= 1'b0;
      compareStage_controlPipe_translated_s2mPipe_rValid <= 1'b0;
      diffStage_mainOnePixelStream_rValid <= 1'b0;
      diffStage_mainOnePixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_counterOnePixelStream_rValid <= 1'b0;
      diffStage_counterOnePixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_mainTwoPixelStream_rValid <= 1'b0;
      diffStage_mainTwoPixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_counterTwoPixelStream_rValid <= 1'b0;
      diffStage_counterTwoPixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_mainThreePixelStream_rValid <= 1'b0;
      diffStage_mainThreePixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_counterThreePixelStream_rValid <= 1'b0;
      diffStage_counterThreePixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_mainOneValidStream_rValid <= 1'b0;
      diffStage_mainOneValidStream_s2mPipe_rValid <= 1'b0;
      diffStage_counterOneValidStream_rValid <= 1'b0;
      diffStage_counterOneValidStream_s2mPipe_rValid <= 1'b0;
      diffStage_mainTwoValidStream_rValid <= 1'b0;
      diffStage_mainTwoValidStream_s2mPipe_rValid <= 1'b0;
      diffStage_counterTwoValidStream_rValid <= 1'b0;
      diffStage_counterTwoValidStream_s2mPipe_rValid <= 1'b0;
      diffStage_mainThreeValidStream_rValid <= 1'b0;
      diffStage_mainThreeValidStream_s2mPipe_rValid <= 1'b0;
      diffStage_counterThreeValidStream_rValid <= 1'b0;
      diffStage_counterThreeValidStream_s2mPipe_rValid <= 1'b0;
      resultStage_controlPipeBeforePipe_rValid <= 1'b0;
      resultStage_controlPipeBeforePipe_s2mPipe_rValid <= 1'b0;
      resultStage_pixelStream_rValid <= 1'b0;
      resultStage_pixelStream_s2mPipe_rValid <= 1'b0;
      pixelsStream_rValid <= 1'b0;
      pixelsStream_s2mPipe_rValid <= 1'b0;
      controlStateMachine_stateReg <= controlStateMachine_enumDef_5_BOOT;
    end else begin
      if(when_SuperResolutionPart3_l72) begin
        inpThreeDone <= 1'b0;
      end
      if(when_SuperResolutionPart3_l75) begin
        readDone <= 1'b0;
      end
      if(when_SuperResolutionPart3_l78) begin
        startRead <= 1'b1;
      end
      if(when_SuperResolutionPart3_l78_1) begin
        startRead <= 1'b0;
      end
      inpThreshold <= thresholdIn;
      bmpWidth <= widthIn;
      bmpHeight <= heightIn;
      if(when_SuperResolutionPart3_l93) begin
        holdBuffer <= 1'b0;
      end
      if(when_SuperResolutionPart3_l96) begin
        writeDone <= 1'b0;
      end
      bufferRowCount_value <= bufferRowCount_valueNext;
      if(when_SuperResolutionPart3_l102) begin
        bufferEnable <= 1'b1;
      end
      if(when_SuperResolutionPart3_l102_1) begin
        bufferEnable <= 1'b0;
      end
      if(inpThreeDone) begin
        bufferReuse <= 1'b0;
      end
      bufferWAddr_value <= bufferWAddr_valueNext;
      outPixelAddr_value <= outPixelAddr_valueNext;
      outRowCount_value <= outRowCount_valueNext;
      alreadySendRow_value <= alreadySendRow_valueNext;
      alreadySendCountInRow_value <= alreadySendCountInRow_valueNext;
      if(when_SuperResolutionPart3_l154) begin
        bufferSwitch <= 2'b00;
        nextRowBuffer <= {1'd0, CICC1851_nextRowBuffer};
        currentRowBuffer <= 2'b00;
        minDiff <= 8'h0;
        candidatePixel <= 8'h0;
        isHorizontalDirection <= 1'b0;
      end
      if(pixelsIn_valid) begin
        pixelsIn_rValid <= 1'b1;
      end
      if(pixelsIn_s2mPipe_ready) begin
        pixelsIn_rValid <= 1'b0;
      end
      if(pixelsIn_s2mPipe_ready) begin
        pixelsIn_s2mPipe_rValid <= pixelsIn_s2mPipe_valid;
      end
      if(when_SuperResolutionPart3_l226) begin
        bufferReachRowEnd <= 1'b1;
      end
      if(when_SuperResolutionPart3_l227) begin
        bufferReachFinalRow <= 1'b1;
      end
      if(when_SuperResolutionPart3_l230) begin
        if(bufferReachFinalRow) begin
          bufferReuse <= 1'b1;
          bufferReachRowEnd <= 1'b0;
          bufferReachFinalRow <= 1'b0;
        end else begin
          bufferReachRowEnd <= 1'b0;
        end
      end
      if(when_SuperResolutionPart3_l243) begin
        if(when_SuperResolutionPart3_l244) begin
          bufferSwitch <= 2'b00;
        end else begin
          bufferSwitch <= (bufferSwitch + 2'b01);
        end
      end
      if(when_SuperResolutionPart3_l251) begin
        holdBuffer <= 1'b1;
        bufferEnable <= 1'b0;
        if(when_SuperResolutionPart3_l255) begin
          writeDone <= 1'b1;
          bufferEnable <= 1'b0;
        end
      end
      if(when_SuperResolutionPart3_l262) begin
        frameStart <= 1'b1;
      end
      if(inpThreeDone) begin
        inpThreeDone <= 1'b0;
      end
      if(when_SuperResolutionPart3_l270) begin
        alreadyReachRowEnd <= 1'b1;
      end
      if(when_SuperResolutionPart3_l271) begin
        alreadyReachFinalRow <= 1'b1;
      end
      if(pixelsOut_fire_2) begin
        if(alreadyReachRowEnd) begin
          alreadyReachRowEnd <= 1'b0;
          if(alreadyReachFinalRow) begin
            alreadyReachFinalRow <= 1'b0;
          end
        end
      end
      if(when_SuperResolutionPart3_l282) begin
        inpThreeDone <= 1'b1;
      end
      if(mainPixelAddrOneStream_valid) begin
        mainPixelAddrOneStream_rValid <= 1'b1;
      end
      if(mainPixelAddrOneStream_s2mPipe_ready) begin
        mainPixelAddrOneStream_rValid <= 1'b0;
      end
      if(mainPixelAddrOneStream_s2mPipe_ready) begin
        mainPixelAddrOneStream_s2mPipe_rValid <= mainPixelAddrOneStream_s2mPipe_valid;
      end
      if(CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(mainPixelAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_2 <= mainPixelAddrOneStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_1) begin
        CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_1) begin
        CICC1851_readStage_mainOnePixelStream_valid <= (CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready || CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_3);
      end
      if(counterPixelAddrOneStream_valid) begin
        counterPixelAddrOneStream_rValid <= 1'b1;
      end
      if(counterPixelAddrOneStream_s2mPipe_ready) begin
        counterPixelAddrOneStream_rValid <= 1'b0;
      end
      if(counterPixelAddrOneStream_s2mPipe_ready) begin
        counterPixelAddrOneStream_s2mPipe_rValid <= counterPixelAddrOneStream_s2mPipe_valid;
      end
      if(CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(counterPixelAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_2 <= counterPixelAddrOneStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_2) begin
        CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_2) begin
        CICC1851_readStage_counterOnePixelStream_valid <= (CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready || CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_3);
      end
      if(mainPixelAddrTwoStream_valid) begin
        mainPixelAddrTwoStream_rValid <= 1'b1;
      end
      if(mainPixelAddrTwoStream_s2mPipe_ready) begin
        mainPixelAddrTwoStream_rValid <= 1'b0;
      end
      if(mainPixelAddrTwoStream_s2mPipe_ready) begin
        mainPixelAddrTwoStream_s2mPipe_rValid <= mainPixelAddrTwoStream_s2mPipe_valid;
      end
      if(CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= mainPixelAddrTwoStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_3) begin
        CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_3) begin
        CICC1851_readStage_mainTwoPixelStream_valid <= (CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready || CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_3);
      end
      if(counterPixelAddrTwoStream_valid) begin
        counterPixelAddrTwoStream_rValid <= 1'b1;
      end
      if(counterPixelAddrTwoStream_s2mPipe_ready) begin
        counterPixelAddrTwoStream_rValid <= 1'b0;
      end
      if(counterPixelAddrTwoStream_s2mPipe_ready) begin
        counterPixelAddrTwoStream_s2mPipe_rValid <= counterPixelAddrTwoStream_s2mPipe_valid;
      end
      if(CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= counterPixelAddrTwoStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_4) begin
        CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_4) begin
        CICC1851_readStage_counterTwoPixelStream_valid <= (CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready || CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_3);
      end
      if(mainPixelAddrThreeStream_valid) begin
        mainPixelAddrThreeStream_rValid <= 1'b1;
      end
      if(mainPixelAddrThreeStream_s2mPipe_ready) begin
        mainPixelAddrThreeStream_rValid <= 1'b0;
      end
      if(mainPixelAddrThreeStream_s2mPipe_ready) begin
        mainPixelAddrThreeStream_s2mPipe_rValid <= mainPixelAddrThreeStream_s2mPipe_valid;
      end
      if(CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_2 <= mainPixelAddrThreeStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_5) begin
        CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_5) begin
        CICC1851_readStage_mainThreePixelStream_valid <= (CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready || CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_3);
      end
      if(counterPixelAddrThreeStream_valid) begin
        counterPixelAddrThreeStream_rValid <= 1'b1;
      end
      if(counterPixelAddrThreeStream_s2mPipe_ready) begin
        counterPixelAddrThreeStream_rValid <= 1'b0;
      end
      if(counterPixelAddrThreeStream_s2mPipe_ready) begin
        counterPixelAddrThreeStream_s2mPipe_rValid <= counterPixelAddrThreeStream_s2mPipe_valid;
      end
      if(CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_2 <= counterPixelAddrThreeStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_6) begin
        CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_6) begin
        CICC1851_readStage_counterThreePixelStream_valid <= (CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready || CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_3);
      end
      if(mainValidAddrOneStream_valid) begin
        mainValidAddrOneStream_rValid <= 1'b1;
      end
      if(mainValidAddrOneStream_s2mPipe_ready) begin
        mainValidAddrOneStream_rValid <= 1'b0;
      end
      if(mainValidAddrOneStream_s2mPipe_ready) begin
        mainValidAddrOneStream_s2mPipe_rValid <= mainValidAddrOneStream_s2mPipe_valid;
      end
      if(CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(mainValidAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_2 <= mainValidAddrOneStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_7) begin
        CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_7) begin
        CICC1851_readStage_mainOneValidStream_valid <= (CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready || CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_3);
      end
      if(counterValidAddrOneStream_valid) begin
        counterValidAddrOneStream_rValid <= 1'b1;
      end
      if(counterValidAddrOneStream_s2mPipe_ready) begin
        counterValidAddrOneStream_rValid <= 1'b0;
      end
      if(counterValidAddrOneStream_s2mPipe_ready) begin
        counterValidAddrOneStream_s2mPipe_rValid <= counterValidAddrOneStream_s2mPipe_valid;
      end
      if(CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(counterValidAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_2 <= counterValidAddrOneStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_8) begin
        CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_8) begin
        CICC1851_readStage_counterOneValidStream_valid <= (CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready || CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_3);
      end
      if(mainValidAddrTwoStream_valid) begin
        mainValidAddrTwoStream_rValid <= 1'b1;
      end
      if(mainValidAddrTwoStream_s2mPipe_ready) begin
        mainValidAddrTwoStream_rValid <= 1'b0;
      end
      if(mainValidAddrTwoStream_s2mPipe_ready) begin
        mainValidAddrTwoStream_s2mPipe_rValid <= mainValidAddrTwoStream_s2mPipe_valid;
      end
      if(CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(mainValidAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= mainValidAddrTwoStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_9) begin
        CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_9) begin
        CICC1851_readStage_mainTwoValidStream_valid <= (CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready || CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_3);
      end
      if(counterValidAddrTwoStream_valid) begin
        counterValidAddrTwoStream_rValid <= 1'b1;
      end
      if(counterValidAddrTwoStream_s2mPipe_ready) begin
        counterValidAddrTwoStream_rValid <= 1'b0;
      end
      if(counterValidAddrTwoStream_s2mPipe_ready) begin
        counterValidAddrTwoStream_s2mPipe_rValid <= counterValidAddrTwoStream_s2mPipe_valid;
      end
      if(CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(counterValidAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= counterValidAddrTwoStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_10) begin
        CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_10) begin
        CICC1851_readStage_counterTwoValidStream_valid <= (CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready || CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_3);
      end
      if(mainValidAddrThreeStream_valid) begin
        mainValidAddrThreeStream_rValid <= 1'b1;
      end
      if(mainValidAddrThreeStream_s2mPipe_ready) begin
        mainValidAddrThreeStream_rValid <= 1'b0;
      end
      if(mainValidAddrThreeStream_s2mPipe_ready) begin
        mainValidAddrThreeStream_s2mPipe_rValid <= mainValidAddrThreeStream_s2mPipe_valid;
      end
      if(CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(mainValidAddrThreeStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_2 <= mainValidAddrThreeStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_11) begin
        CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_11) begin
        CICC1851_readStage_mainThreeValidStream_valid <= (CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready || CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_3);
      end
      if(counterValidAddrThreeStream_valid) begin
        counterValidAddrThreeStream_rValid <= 1'b1;
      end
      if(counterValidAddrThreeStream_s2mPipe_ready) begin
        counterValidAddrThreeStream_rValid <= 1'b0;
      end
      if(counterValidAddrThreeStream_s2mPipe_ready) begin
        counterValidAddrThreeStream_s2mPipe_rValid <= counterValidAddrThreeStream_s2mPipe_valid;
      end
      if(CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(counterValidAddrThreeStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_2 <= counterValidAddrThreeStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_12) begin
        CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_12) begin
        CICC1851_readStage_counterThreeValidStream_valid <= (CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready || CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_3);
      end
      if(controlStream_valid) begin
        controlStream_rValid <= 1'b1;
      end
      if(controlStream_s2mPipe_ready) begin
        controlStream_rValid <= 1'b0;
      end
      if(controlStream_s2mPipe_ready) begin
        controlStream_s2mPipe_rValid <= controlStream_s2mPipe_valid;
      end
      if(controlStream_s2mPipe_m2sPipe_ready) begin
        controlStream_s2mPipe_m2sPipe_rValid <= controlStream_s2mPipe_m2sPipe_valid;
      end
      if(controlStream_s2mPipe_m2sPipe_m2sPipe_valid) begin
        controlStream_s2mPipe_m2sPipe_m2sPipe_rValid <= 1'b1;
      end
      if(controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready) begin
        controlStream_s2mPipe_m2sPipe_m2sPipe_rValid <= 1'b0;
      end
      if(controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready) begin
        controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_valid;
      end
      if(readStage_mainOnePixelStream_valid) begin
        readStage_mainOnePixelStream_rValid <= 1'b1;
      end
      if(readStage_mainOnePixelStream_s2mPipe_ready) begin
        readStage_mainOnePixelStream_rValid <= 1'b0;
      end
      if(readStage_mainOnePixelStream_s2mPipe_ready) begin
        readStage_mainOnePixelStream_s2mPipe_rValid <= readStage_mainOnePixelStream_s2mPipe_valid;
      end
      if(readStage_counterOnePixelStream_valid) begin
        readStage_counterOnePixelStream_rValid <= 1'b1;
      end
      if(readStage_counterOnePixelStream_s2mPipe_ready) begin
        readStage_counterOnePixelStream_rValid <= 1'b0;
      end
      if(readStage_counterOnePixelStream_s2mPipe_ready) begin
        readStage_counterOnePixelStream_s2mPipe_rValid <= readStage_counterOnePixelStream_s2mPipe_valid;
      end
      if(readStage_mainTwoPixelStream_valid) begin
        readStage_mainTwoPixelStream_rValid <= 1'b1;
      end
      if(readStage_mainTwoPixelStream_s2mPipe_ready) begin
        readStage_mainTwoPixelStream_rValid <= 1'b0;
      end
      if(readStage_mainTwoPixelStream_s2mPipe_ready) begin
        readStage_mainTwoPixelStream_s2mPipe_rValid <= readStage_mainTwoPixelStream_s2mPipe_valid;
      end
      if(readStage_counterTwoPixelStream_valid) begin
        readStage_counterTwoPixelStream_rValid <= 1'b1;
      end
      if(readStage_counterTwoPixelStream_s2mPipe_ready) begin
        readStage_counterTwoPixelStream_rValid <= 1'b0;
      end
      if(readStage_counterTwoPixelStream_s2mPipe_ready) begin
        readStage_counterTwoPixelStream_s2mPipe_rValid <= readStage_counterTwoPixelStream_s2mPipe_valid;
      end
      if(readStage_mainThreePixelStream_valid) begin
        readStage_mainThreePixelStream_rValid <= 1'b1;
      end
      if(readStage_mainThreePixelStream_s2mPipe_ready) begin
        readStage_mainThreePixelStream_rValid <= 1'b0;
      end
      if(readStage_mainThreePixelStream_s2mPipe_ready) begin
        readStage_mainThreePixelStream_s2mPipe_rValid <= readStage_mainThreePixelStream_s2mPipe_valid;
      end
      if(readStage_counterThreePixelStream_valid) begin
        readStage_counterThreePixelStream_rValid <= 1'b1;
      end
      if(readStage_counterThreePixelStream_s2mPipe_ready) begin
        readStage_counterThreePixelStream_rValid <= 1'b0;
      end
      if(readStage_counterThreePixelStream_s2mPipe_ready) begin
        readStage_counterThreePixelStream_s2mPipe_rValid <= readStage_counterThreePixelStream_s2mPipe_valid;
      end
      if(readStage_mainOneValidStream_valid) begin
        readStage_mainOneValidStream_rValid <= 1'b1;
      end
      if(readStage_mainOneValidStream_s2mPipe_ready) begin
        readStage_mainOneValidStream_rValid <= 1'b0;
      end
      if(readStage_mainOneValidStream_s2mPipe_ready) begin
        readStage_mainOneValidStream_s2mPipe_rValid <= readStage_mainOneValidStream_s2mPipe_valid;
      end
      if(readStage_counterOneValidStream_valid) begin
        readStage_counterOneValidStream_rValid <= 1'b1;
      end
      if(readStage_counterOneValidStream_s2mPipe_ready) begin
        readStage_counterOneValidStream_rValid <= 1'b0;
      end
      if(readStage_counterOneValidStream_s2mPipe_ready) begin
        readStage_counterOneValidStream_s2mPipe_rValid <= readStage_counterOneValidStream_s2mPipe_valid;
      end
      if(readStage_mainTwoValidStream_valid) begin
        readStage_mainTwoValidStream_rValid <= 1'b1;
      end
      if(readStage_mainTwoValidStream_s2mPipe_ready) begin
        readStage_mainTwoValidStream_rValid <= 1'b0;
      end
      if(readStage_mainTwoValidStream_s2mPipe_ready) begin
        readStage_mainTwoValidStream_s2mPipe_rValid <= readStage_mainTwoValidStream_s2mPipe_valid;
      end
      if(readStage_counterTwoValidStream_valid) begin
        readStage_counterTwoValidStream_rValid <= 1'b1;
      end
      if(readStage_counterTwoValidStream_s2mPipe_ready) begin
        readStage_counterTwoValidStream_rValid <= 1'b0;
      end
      if(readStage_counterTwoValidStream_s2mPipe_ready) begin
        readStage_counterTwoValidStream_s2mPipe_rValid <= readStage_counterTwoValidStream_s2mPipe_valid;
      end
      if(readStage_mainThreeValidStream_valid) begin
        readStage_mainThreeValidStream_rValid <= 1'b1;
      end
      if(readStage_mainThreeValidStream_s2mPipe_ready) begin
        readStage_mainThreeValidStream_rValid <= 1'b0;
      end
      if(readStage_mainThreeValidStream_s2mPipe_ready) begin
        readStage_mainThreeValidStream_s2mPipe_rValid <= readStage_mainThreeValidStream_s2mPipe_valid;
      end
      if(readStage_counterThreeValidStream_valid) begin
        readStage_counterThreeValidStream_rValid <= 1'b1;
      end
      if(readStage_counterThreeValidStream_s2mPipe_ready) begin
        readStage_counterThreeValidStream_rValid <= 1'b0;
      end
      if(readStage_counterThreeValidStream_s2mPipe_ready) begin
        readStage_counterThreeValidStream_s2mPipe_rValid <= readStage_counterThreeValidStream_s2mPipe_valid;
      end
      if(readStage_controlPipe_translated_valid) begin
        readStage_controlPipe_translated_rValid <= 1'b1;
      end
      if(readStage_controlPipe_translated_s2mPipe_ready) begin
        readStage_controlPipe_translated_rValid <= 1'b0;
      end
      if(readStage_controlPipe_translated_s2mPipe_ready) begin
        readStage_controlPipe_translated_s2mPipe_rValid <= readStage_controlPipe_translated_s2mPipe_valid;
      end
      if(compareStage_mainOnePixelStream_valid) begin
        compareStage_mainOnePixelStream_rValid <= 1'b1;
      end
      if(compareStage_mainOnePixelStream_s2mPipe_ready) begin
        compareStage_mainOnePixelStream_rValid <= 1'b0;
      end
      if(compareStage_mainOnePixelStream_s2mPipe_ready) begin
        compareStage_mainOnePixelStream_s2mPipe_rValid <= compareStage_mainOnePixelStream_s2mPipe_valid;
      end
      if(compareStage_counterOnePixelStream_valid) begin
        compareStage_counterOnePixelStream_rValid <= 1'b1;
      end
      if(compareStage_counterOnePixelStream_s2mPipe_ready) begin
        compareStage_counterOnePixelStream_rValid <= 1'b0;
      end
      if(compareStage_counterOnePixelStream_s2mPipe_ready) begin
        compareStage_counterOnePixelStream_s2mPipe_rValid <= compareStage_counterOnePixelStream_s2mPipe_valid;
      end
      if(compareStage_mainTwoPixelStream_valid) begin
        compareStage_mainTwoPixelStream_rValid <= 1'b1;
      end
      if(compareStage_mainTwoPixelStream_s2mPipe_ready) begin
        compareStage_mainTwoPixelStream_rValid <= 1'b0;
      end
      if(compareStage_mainTwoPixelStream_s2mPipe_ready) begin
        compareStage_mainTwoPixelStream_s2mPipe_rValid <= compareStage_mainTwoPixelStream_s2mPipe_valid;
      end
      if(compareStage_counterTwoPixelStream_valid) begin
        compareStage_counterTwoPixelStream_rValid <= 1'b1;
      end
      if(compareStage_counterTwoPixelStream_s2mPipe_ready) begin
        compareStage_counterTwoPixelStream_rValid <= 1'b0;
      end
      if(compareStage_counterTwoPixelStream_s2mPipe_ready) begin
        compareStage_counterTwoPixelStream_s2mPipe_rValid <= compareStage_counterTwoPixelStream_s2mPipe_valid;
      end
      if(compareStage_mainThreePixelStream_valid) begin
        compareStage_mainThreePixelStream_rValid <= 1'b1;
      end
      if(compareStage_mainThreePixelStream_s2mPipe_ready) begin
        compareStage_mainThreePixelStream_rValid <= 1'b0;
      end
      if(compareStage_mainThreePixelStream_s2mPipe_ready) begin
        compareStage_mainThreePixelStream_s2mPipe_rValid <= compareStage_mainThreePixelStream_s2mPipe_valid;
      end
      if(compareStage_counterThreePixelStream_valid) begin
        compareStage_counterThreePixelStream_rValid <= 1'b1;
      end
      if(compareStage_counterThreePixelStream_s2mPipe_ready) begin
        compareStage_counterThreePixelStream_rValid <= 1'b0;
      end
      if(compareStage_counterThreePixelStream_s2mPipe_ready) begin
        compareStage_counterThreePixelStream_s2mPipe_rValid <= compareStage_counterThreePixelStream_s2mPipe_valid;
      end
      if(compareStage_mainOneValidStream_valid) begin
        compareStage_mainOneValidStream_rValid <= 1'b1;
      end
      if(compareStage_mainOneValidStream_s2mPipe_ready) begin
        compareStage_mainOneValidStream_rValid <= 1'b0;
      end
      if(compareStage_mainOneValidStream_s2mPipe_ready) begin
        compareStage_mainOneValidStream_s2mPipe_rValid <= compareStage_mainOneValidStream_s2mPipe_valid;
      end
      if(compareStage_counterOneValidStream_valid) begin
        compareStage_counterOneValidStream_rValid <= 1'b1;
      end
      if(compareStage_counterOneValidStream_s2mPipe_ready) begin
        compareStage_counterOneValidStream_rValid <= 1'b0;
      end
      if(compareStage_counterOneValidStream_s2mPipe_ready) begin
        compareStage_counterOneValidStream_s2mPipe_rValid <= compareStage_counterOneValidStream_s2mPipe_valid;
      end
      if(compareStage_mainTwoValidStream_valid) begin
        compareStage_mainTwoValidStream_rValid <= 1'b1;
      end
      if(compareStage_mainTwoValidStream_s2mPipe_ready) begin
        compareStage_mainTwoValidStream_rValid <= 1'b0;
      end
      if(compareStage_mainTwoValidStream_s2mPipe_ready) begin
        compareStage_mainTwoValidStream_s2mPipe_rValid <= compareStage_mainTwoValidStream_s2mPipe_valid;
      end
      if(compareStage_counterTwoValidStream_valid) begin
        compareStage_counterTwoValidStream_rValid <= 1'b1;
      end
      if(compareStage_counterTwoValidStream_s2mPipe_ready) begin
        compareStage_counterTwoValidStream_rValid <= 1'b0;
      end
      if(compareStage_counterTwoValidStream_s2mPipe_ready) begin
        compareStage_counterTwoValidStream_s2mPipe_rValid <= compareStage_counterTwoValidStream_s2mPipe_valid;
      end
      if(compareStage_mainThreeValidStream_valid) begin
        compareStage_mainThreeValidStream_rValid <= 1'b1;
      end
      if(compareStage_mainThreeValidStream_s2mPipe_ready) begin
        compareStage_mainThreeValidStream_rValid <= 1'b0;
      end
      if(compareStage_mainThreeValidStream_s2mPipe_ready) begin
        compareStage_mainThreeValidStream_s2mPipe_rValid <= compareStage_mainThreeValidStream_s2mPipe_valid;
      end
      if(compareStage_counterThreeValidStream_valid) begin
        compareStage_counterThreeValidStream_rValid <= 1'b1;
      end
      if(compareStage_counterThreeValidStream_s2mPipe_ready) begin
        compareStage_counterThreeValidStream_rValid <= 1'b0;
      end
      if(compareStage_counterThreeValidStream_s2mPipe_ready) begin
        compareStage_counterThreeValidStream_s2mPipe_rValid <= compareStage_counterThreeValidStream_s2mPipe_valid;
      end
      if(compareStage_controlPipe_translated_valid) begin
        compareStage_controlPipe_translated_rValid <= 1'b1;
      end
      if(compareStage_controlPipe_translated_s2mPipe_ready) begin
        compareStage_controlPipe_translated_rValid <= 1'b0;
      end
      if(compareStage_controlPipe_translated_s2mPipe_ready) begin
        compareStage_controlPipe_translated_s2mPipe_rValid <= compareStage_controlPipe_translated_s2mPipe_valid;
      end
      if(diffStage_mainOnePixelStream_valid) begin
        diffStage_mainOnePixelStream_rValid <= 1'b1;
      end
      if(diffStage_mainOnePixelStream_s2mPipe_ready) begin
        diffStage_mainOnePixelStream_rValid <= 1'b0;
      end
      if(diffStage_mainOnePixelStream_s2mPipe_ready) begin
        diffStage_mainOnePixelStream_s2mPipe_rValid <= diffStage_mainOnePixelStream_s2mPipe_valid;
      end
      if(diffStage_counterOnePixelStream_valid) begin
        diffStage_counterOnePixelStream_rValid <= 1'b1;
      end
      if(diffStage_counterOnePixelStream_s2mPipe_ready) begin
        diffStage_counterOnePixelStream_rValid <= 1'b0;
      end
      if(diffStage_counterOnePixelStream_s2mPipe_ready) begin
        diffStage_counterOnePixelStream_s2mPipe_rValid <= diffStage_counterOnePixelStream_s2mPipe_valid;
      end
      if(diffStage_mainTwoPixelStream_valid) begin
        diffStage_mainTwoPixelStream_rValid <= 1'b1;
      end
      if(diffStage_mainTwoPixelStream_s2mPipe_ready) begin
        diffStage_mainTwoPixelStream_rValid <= 1'b0;
      end
      if(diffStage_mainTwoPixelStream_s2mPipe_ready) begin
        diffStage_mainTwoPixelStream_s2mPipe_rValid <= diffStage_mainTwoPixelStream_s2mPipe_valid;
      end
      if(diffStage_counterTwoPixelStream_valid) begin
        diffStage_counterTwoPixelStream_rValid <= 1'b1;
      end
      if(diffStage_counterTwoPixelStream_s2mPipe_ready) begin
        diffStage_counterTwoPixelStream_rValid <= 1'b0;
      end
      if(diffStage_counterTwoPixelStream_s2mPipe_ready) begin
        diffStage_counterTwoPixelStream_s2mPipe_rValid <= diffStage_counterTwoPixelStream_s2mPipe_valid;
      end
      if(diffStage_mainThreePixelStream_valid) begin
        diffStage_mainThreePixelStream_rValid <= 1'b1;
      end
      if(diffStage_mainThreePixelStream_s2mPipe_ready) begin
        diffStage_mainThreePixelStream_rValid <= 1'b0;
      end
      if(diffStage_mainThreePixelStream_s2mPipe_ready) begin
        diffStage_mainThreePixelStream_s2mPipe_rValid <= diffStage_mainThreePixelStream_s2mPipe_valid;
      end
      if(diffStage_counterThreePixelStream_valid) begin
        diffStage_counterThreePixelStream_rValid <= 1'b1;
      end
      if(diffStage_counterThreePixelStream_s2mPipe_ready) begin
        diffStage_counterThreePixelStream_rValid <= 1'b0;
      end
      if(diffStage_counterThreePixelStream_s2mPipe_ready) begin
        diffStage_counterThreePixelStream_s2mPipe_rValid <= diffStage_counterThreePixelStream_s2mPipe_valid;
      end
      if(diffStage_mainOneValidStream_valid) begin
        diffStage_mainOneValidStream_rValid <= 1'b1;
      end
      if(diffStage_mainOneValidStream_s2mPipe_ready) begin
        diffStage_mainOneValidStream_rValid <= 1'b0;
      end
      if(diffStage_mainOneValidStream_s2mPipe_ready) begin
        diffStage_mainOneValidStream_s2mPipe_rValid <= diffStage_mainOneValidStream_s2mPipe_valid;
      end
      if(diffStage_counterOneValidStream_valid) begin
        diffStage_counterOneValidStream_rValid <= 1'b1;
      end
      if(diffStage_counterOneValidStream_s2mPipe_ready) begin
        diffStage_counterOneValidStream_rValid <= 1'b0;
      end
      if(diffStage_counterOneValidStream_s2mPipe_ready) begin
        diffStage_counterOneValidStream_s2mPipe_rValid <= diffStage_counterOneValidStream_s2mPipe_valid;
      end
      if(diffStage_mainTwoValidStream_valid) begin
        diffStage_mainTwoValidStream_rValid <= 1'b1;
      end
      if(diffStage_mainTwoValidStream_s2mPipe_ready) begin
        diffStage_mainTwoValidStream_rValid <= 1'b0;
      end
      if(diffStage_mainTwoValidStream_s2mPipe_ready) begin
        diffStage_mainTwoValidStream_s2mPipe_rValid <= diffStage_mainTwoValidStream_s2mPipe_valid;
      end
      if(diffStage_counterTwoValidStream_valid) begin
        diffStage_counterTwoValidStream_rValid <= 1'b1;
      end
      if(diffStage_counterTwoValidStream_s2mPipe_ready) begin
        diffStage_counterTwoValidStream_rValid <= 1'b0;
      end
      if(diffStage_counterTwoValidStream_s2mPipe_ready) begin
        diffStage_counterTwoValidStream_s2mPipe_rValid <= diffStage_counterTwoValidStream_s2mPipe_valid;
      end
      if(diffStage_mainThreeValidStream_valid) begin
        diffStage_mainThreeValidStream_rValid <= 1'b1;
      end
      if(diffStage_mainThreeValidStream_s2mPipe_ready) begin
        diffStage_mainThreeValidStream_rValid <= 1'b0;
      end
      if(diffStage_mainThreeValidStream_s2mPipe_ready) begin
        diffStage_mainThreeValidStream_s2mPipe_rValid <= diffStage_mainThreeValidStream_s2mPipe_valid;
      end
      if(diffStage_counterThreeValidStream_valid) begin
        diffStage_counterThreeValidStream_rValid <= 1'b1;
      end
      if(diffStage_counterThreeValidStream_s2mPipe_ready) begin
        diffStage_counterThreeValidStream_rValid <= 1'b0;
      end
      if(diffStage_counterThreeValidStream_s2mPipe_ready) begin
        diffStage_counterThreeValidStream_s2mPipe_rValid <= diffStage_counterThreeValidStream_s2mPipe_valid;
      end
      if(resultStage_controlPipeBeforePipe_valid) begin
        resultStage_controlPipeBeforePipe_rValid <= 1'b1;
      end
      if(resultStage_controlPipeBeforePipe_s2mPipe_ready) begin
        resultStage_controlPipeBeforePipe_rValid <= 1'b0;
      end
      if(resultStage_controlPipeBeforePipe_s2mPipe_ready) begin
        resultStage_controlPipeBeforePipe_s2mPipe_rValid <= resultStage_controlPipeBeforePipe_s2mPipe_valid;
      end
      if(resultStage_pixelStream_valid) begin
        resultStage_pixelStream_rValid <= 1'b1;
      end
      if(resultStage_pixelStream_s2mPipe_ready) begin
        resultStage_pixelStream_rValid <= 1'b0;
      end
      if(resultStage_pixelStream_s2mPipe_ready) begin
        resultStage_pixelStream_s2mPipe_rValid <= resultStage_pixelStream_s2mPipe_valid;
      end
      if(when_SuperResolutionPart3_l1115) begin
        isHorizontalDirection <= resultStage_controlPipeBeforePipe_payload_isHorizontalMin;
        minDiff <= resultStage_controlPipeBeforePipe_payload_minDiff;
        candidatePixel <= resultStage_pixelStream_payload;
      end
      if(diffStage_controlPipe_fire) begin
        inValidMinDiff <= diffStage_controlPipe_payload_inValidMinDiff;
      end
      if(pixelsStream_valid) begin
        pixelsStream_rValid <= 1'b1;
      end
      if(pixelsStream_s2mPipe_ready) begin
        pixelsStream_rValid <= 1'b0;
      end
      if(pixelsStream_s2mPipe_ready) begin
        pixelsStream_s2mPipe_rValid <= pixelsStream_s2mPipe_valid;
      end
      controlStateMachine_stateReg <= controlStateMachine_stateNext;
      case(controlStateMachine_stateReg)
        controlStateMachine_enumDef_5_HOLD : begin
        end
        controlStateMachine_enumDef_5_PASS : begin
        end
        controlStateMachine_enumDef_5_EXTRA : begin
          if(when_SuperResolutionPart3_l1220) begin
            frameStart <= 1'b0;
          end
          if(when_SuperResolutionPart3_l1223) begin
            outReachRowEnd <= 1'b1;
          end
          if(when_SuperResolutionPart3_l1224) begin
            outReachFinalRow <= 1'b1;
          end
          if(when_SuperResolutionPart3_l1226) begin
            if(outReachFinalRow) begin
              startRead <= 1'b0;
              readDone <= 1'b1;
              outReachRowEnd <= 1'b0;
              outReachFinalRow <= 1'b0;
            end else begin
              outReachRowEnd <= 1'b0;
            end
          end
          if(controlStream_fire_6) begin
            if(outReachRowEnd) begin
              outReachRowEnd <= 1'b0;
            end
          end
          if(when_SuperResolutionPart3_l1247) begin
            if(when_SuperResolutionPart3_l1248) begin
              holdBuffer <= 1'b0;
            end
            if(when_SuperResolutionPart3_l1250) begin
              currentRowBuffer <= 2'b00;
            end else begin
              currentRowBuffer <= (currentRowBuffer + 2'b01);
            end
            if(when_SuperResolutionPart3_l1252) begin
              nextRowBuffer <= 2'b00;
            end else begin
              nextRowBuffer <= (nextRowBuffer + 2'b01);
            end
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(posedge clk) begin
    startIn_regNext <= startIn;
    startIn_regNext_1 <= startIn;
    if(pixelsIn_ready) begin
      pixelsIn_rData_pixel <= pixelsIn_payload_pixel;
      pixelsIn_rData_frameStart <= pixelsIn_payload_frameStart;
      pixelsIn_rData_rowEnd <= pixelsIn_payload_rowEnd;
      pixelsIn_rData_inpValid <= pixelsIn_payload_inpValid;
    end
    if(pixelsIn_s2mPipe_ready) begin
      pixelsIn_s2mPipe_rData_pixel <= pixelsIn_s2mPipe_payload_pixel;
      pixelsIn_s2mPipe_rData_frameStart <= pixelsIn_s2mPipe_payload_frameStart;
      pixelsIn_s2mPipe_rData_rowEnd <= pixelsIn_s2mPipe_payload_rowEnd;
      pixelsIn_s2mPipe_rData_inpValid <= pixelsIn_s2mPipe_payload_inpValid;
    end
    if(mainPixelAddrOneStream_ready) begin
      mainPixelAddrOneStream_rData <= mainPixelAddrOneStream_payload;
    end
    if(mainPixelAddrOneStream_s2mPipe_ready) begin
      mainPixelAddrOneStream_s2mPipe_rData <= mainPixelAddrOneStream_s2mPipe_payload;
    end
    if(CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_mainOnePixelStream_payload_1 <= CICC1851_readStage_mainOnePixelStream_payload;
    end
    if(CICC1851_1) begin
      CICC1851_readStage_mainOnePixelStream_payload_2 <= (CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_mainOnePixelStream_payload_1 : CICC1851_readStage_mainOnePixelStream_payload);
    end
    if(counterPixelAddrOneStream_ready) begin
      counterPixelAddrOneStream_rData <= counterPixelAddrOneStream_payload;
    end
    if(counterPixelAddrOneStream_s2mPipe_ready) begin
      counterPixelAddrOneStream_s2mPipe_rData <= counterPixelAddrOneStream_s2mPipe_payload;
    end
    if(CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_counterOnePixelStream_payload_1 <= CICC1851_readStage_counterOnePixelStream_payload;
    end
    if(CICC1851_2) begin
      CICC1851_readStage_counterOnePixelStream_payload_2 <= (CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_counterOnePixelStream_payload_1 : CICC1851_readStage_counterOnePixelStream_payload);
    end
    if(mainPixelAddrTwoStream_ready) begin
      mainPixelAddrTwoStream_rData <= mainPixelAddrTwoStream_payload;
    end
    if(mainPixelAddrTwoStream_s2mPipe_ready) begin
      mainPixelAddrTwoStream_s2mPipe_rData <= mainPixelAddrTwoStream_s2mPipe_payload;
    end
    if(CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_mainTwoPixelStream_payload_1 <= CICC1851_readStage_mainTwoPixelStream_payload;
    end
    if(CICC1851_3) begin
      CICC1851_readStage_mainTwoPixelStream_payload_2 <= (CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_mainTwoPixelStream_payload_1 : CICC1851_readStage_mainTwoPixelStream_payload);
    end
    if(counterPixelAddrTwoStream_ready) begin
      counterPixelAddrTwoStream_rData <= counterPixelAddrTwoStream_payload;
    end
    if(counterPixelAddrTwoStream_s2mPipe_ready) begin
      counterPixelAddrTwoStream_s2mPipe_rData <= counterPixelAddrTwoStream_s2mPipe_payload;
    end
    if(CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_counterTwoPixelStream_payload_1 <= CICC1851_readStage_counterTwoPixelStream_payload;
    end
    if(CICC1851_4) begin
      CICC1851_readStage_counterTwoPixelStream_payload_2 <= (CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_counterTwoPixelStream_payload_1 : CICC1851_readStage_counterTwoPixelStream_payload);
    end
    if(mainPixelAddrThreeStream_ready) begin
      mainPixelAddrThreeStream_rData <= mainPixelAddrThreeStream_payload;
    end
    if(mainPixelAddrThreeStream_s2mPipe_ready) begin
      mainPixelAddrThreeStream_s2mPipe_rData <= mainPixelAddrThreeStream_s2mPipe_payload;
    end
    if(CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_mainThreePixelStream_payload_1 <= CICC1851_readStage_mainThreePixelStream_payload;
    end
    if(CICC1851_5) begin
      CICC1851_readStage_mainThreePixelStream_payload_2 <= (CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_mainThreePixelStream_payload_1 : CICC1851_readStage_mainThreePixelStream_payload);
    end
    if(counterPixelAddrThreeStream_ready) begin
      counterPixelAddrThreeStream_rData <= counterPixelAddrThreeStream_payload;
    end
    if(counterPixelAddrThreeStream_s2mPipe_ready) begin
      counterPixelAddrThreeStream_s2mPipe_rData <= counterPixelAddrThreeStream_s2mPipe_payload;
    end
    if(CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_counterThreePixelStream_payload_1 <= CICC1851_readStage_counterThreePixelStream_payload;
    end
    if(CICC1851_6) begin
      CICC1851_readStage_counterThreePixelStream_payload_2 <= (CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_counterThreePixelStream_payload_1 : CICC1851_readStage_counterThreePixelStream_payload);
    end
    if(mainValidAddrOneStream_ready) begin
      mainValidAddrOneStream_rData <= mainValidAddrOneStream_payload;
    end
    if(mainValidAddrOneStream_s2mPipe_ready) begin
      mainValidAddrOneStream_s2mPipe_rData <= mainValidAddrOneStream_s2mPipe_payload;
    end
    if(CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_mainOneValidStream_payload_1 <= CICC1851_readStage_mainOneValidStream_payload;
    end
    if(CICC1851_7) begin
      CICC1851_readStage_mainOneValidStream_payload_2 <= (CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_mainOneValidStream_payload_1 : CICC1851_readStage_mainOneValidStream_payload);
    end
    if(counterValidAddrOneStream_ready) begin
      counterValidAddrOneStream_rData <= counterValidAddrOneStream_payload;
    end
    if(counterValidAddrOneStream_s2mPipe_ready) begin
      counterValidAddrOneStream_s2mPipe_rData <= counterValidAddrOneStream_s2mPipe_payload;
    end
    if(CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_counterOneValidStream_payload_1 <= CICC1851_readStage_counterOneValidStream_payload;
    end
    if(CICC1851_8) begin
      CICC1851_readStage_counterOneValidStream_payload_2 <= (CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_counterOneValidStream_payload_1 : CICC1851_readStage_counterOneValidStream_payload);
    end
    if(mainValidAddrTwoStream_ready) begin
      mainValidAddrTwoStream_rData <= mainValidAddrTwoStream_payload;
    end
    if(mainValidAddrTwoStream_s2mPipe_ready) begin
      mainValidAddrTwoStream_s2mPipe_rData <= mainValidAddrTwoStream_s2mPipe_payload;
    end
    if(CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_mainTwoValidStream_payload_1 <= CICC1851_readStage_mainTwoValidStream_payload;
    end
    if(CICC1851_9) begin
      CICC1851_readStage_mainTwoValidStream_payload_2 <= (CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_mainTwoValidStream_payload_1 : CICC1851_readStage_mainTwoValidStream_payload);
    end
    if(counterValidAddrTwoStream_ready) begin
      counterValidAddrTwoStream_rData <= counterValidAddrTwoStream_payload;
    end
    if(counterValidAddrTwoStream_s2mPipe_ready) begin
      counterValidAddrTwoStream_s2mPipe_rData <= counterValidAddrTwoStream_s2mPipe_payload;
    end
    if(CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_counterTwoValidStream_payload_1 <= CICC1851_readStage_counterTwoValidStream_payload;
    end
    if(CICC1851_10) begin
      CICC1851_readStage_counterTwoValidStream_payload_2 <= (CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_counterTwoValidStream_payload_1 : CICC1851_readStage_counterTwoValidStream_payload);
    end
    if(mainValidAddrThreeStream_ready) begin
      mainValidAddrThreeStream_rData <= mainValidAddrThreeStream_payload;
    end
    if(mainValidAddrThreeStream_s2mPipe_ready) begin
      mainValidAddrThreeStream_s2mPipe_rData <= mainValidAddrThreeStream_s2mPipe_payload;
    end
    if(CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_mainThreeValidStream_payload_1 <= CICC1851_readStage_mainThreeValidStream_payload;
    end
    if(CICC1851_11) begin
      CICC1851_readStage_mainThreeValidStream_payload_2 <= (CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_mainThreeValidStream_payload_1 : CICC1851_readStage_mainThreeValidStream_payload);
    end
    if(counterValidAddrThreeStream_ready) begin
      counterValidAddrThreeStream_rData <= counterValidAddrThreeStream_payload;
    end
    if(counterValidAddrThreeStream_s2mPipe_ready) begin
      counterValidAddrThreeStream_s2mPipe_rData <= counterValidAddrThreeStream_s2mPipe_payload;
    end
    if(CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_counterThreeValidStream_payload_1 <= CICC1851_readStage_counterThreeValidStream_payload;
    end
    if(CICC1851_12) begin
      CICC1851_readStage_counterThreeValidStream_payload_2 <= (CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_counterThreeValidStream_payload_1 : CICC1851_readStage_counterThreeValidStream_payload);
    end
    if(controlStream_ready) begin
      controlStream_rData_frameStart <= controlStream_payload_frameStart;
      controlStream_rData_rowEnd <= controlStream_payload_rowEnd;
      controlStream_rData_pipeValid <= controlStream_payload_pipeValid;
      controlStream_rData_firstRow <= controlStream_payload_firstRow;
      controlStream_rData_lastRow <= controlStream_payload_lastRow;
      controlStream_rData_finalResult <= controlStream_payload_finalResult;
      controlStream_rData_mainCompare <= controlStream_payload_mainCompare;
      controlStream_rData_counterCompare <= controlStream_payload_counterCompare;
      controlStream_rData_horizontalCompare <= controlStream_payload_horizontalCompare;
      controlStream_rData_verticalCompare <= controlStream_payload_verticalCompare;
      controlStream_rData_mainDiff <= controlStream_payload_mainDiff;
      controlStream_rData_counterDiff <= controlStream_payload_counterDiff;
      controlStream_rData_horizontalDiff <= controlStream_payload_horizontalDiff;
      controlStream_rData_verticalDiff <= controlStream_payload_verticalDiff;
      controlStream_rData_isHorizontalMin <= controlStream_payload_isHorizontalMin;
      controlStream_rData_minDiff <= controlStream_payload_minDiff;
      controlStream_rData_currentPosition <= controlStream_payload_currentPosition;
      controlStream_rData_nextPosition <= controlStream_payload_nextPosition;
      controlStream_rData_horizontalDirectionValid <= controlStream_payload_horizontalDirectionValid;
      controlStream_rData_verticalDirectionValid <= controlStream_payload_verticalDirectionValid;
      controlStream_rData_mainDirectionValid <= controlStream_payload_mainDirectionValid;
      controlStream_rData_counterDirectionValid <= controlStream_payload_counterDirectionValid;
      controlStream_rData_inValidMinDiff <= controlStream_payload_inValidMinDiff;
    end
    if(controlStream_s2mPipe_ready) begin
      controlStream_s2mPipe_rData_frameStart <= controlStream_s2mPipe_payload_frameStart;
      controlStream_s2mPipe_rData_rowEnd <= controlStream_s2mPipe_payload_rowEnd;
      controlStream_s2mPipe_rData_pipeValid <= controlStream_s2mPipe_payload_pipeValid;
      controlStream_s2mPipe_rData_firstRow <= controlStream_s2mPipe_payload_firstRow;
      controlStream_s2mPipe_rData_lastRow <= controlStream_s2mPipe_payload_lastRow;
      controlStream_s2mPipe_rData_finalResult <= controlStream_s2mPipe_payload_finalResult;
      controlStream_s2mPipe_rData_mainCompare <= controlStream_s2mPipe_payload_mainCompare;
      controlStream_s2mPipe_rData_counterCompare <= controlStream_s2mPipe_payload_counterCompare;
      controlStream_s2mPipe_rData_horizontalCompare <= controlStream_s2mPipe_payload_horizontalCompare;
      controlStream_s2mPipe_rData_verticalCompare <= controlStream_s2mPipe_payload_verticalCompare;
      controlStream_s2mPipe_rData_mainDiff <= controlStream_s2mPipe_payload_mainDiff;
      controlStream_s2mPipe_rData_counterDiff <= controlStream_s2mPipe_payload_counterDiff;
      controlStream_s2mPipe_rData_horizontalDiff <= controlStream_s2mPipe_payload_horizontalDiff;
      controlStream_s2mPipe_rData_verticalDiff <= controlStream_s2mPipe_payload_verticalDiff;
      controlStream_s2mPipe_rData_isHorizontalMin <= controlStream_s2mPipe_payload_isHorizontalMin;
      controlStream_s2mPipe_rData_minDiff <= controlStream_s2mPipe_payload_minDiff;
      controlStream_s2mPipe_rData_currentPosition <= controlStream_s2mPipe_payload_currentPosition;
      controlStream_s2mPipe_rData_nextPosition <= controlStream_s2mPipe_payload_nextPosition;
      controlStream_s2mPipe_rData_horizontalDirectionValid <= controlStream_s2mPipe_payload_horizontalDirectionValid;
      controlStream_s2mPipe_rData_verticalDirectionValid <= controlStream_s2mPipe_payload_verticalDirectionValid;
      controlStream_s2mPipe_rData_mainDirectionValid <= controlStream_s2mPipe_payload_mainDirectionValid;
      controlStream_s2mPipe_rData_counterDirectionValid <= controlStream_s2mPipe_payload_counterDirectionValid;
      controlStream_s2mPipe_rData_inValidMinDiff <= controlStream_s2mPipe_payload_inValidMinDiff;
    end
    if(controlStream_s2mPipe_m2sPipe_ready) begin
      controlStream_s2mPipe_m2sPipe_rData_frameStart <= controlStream_s2mPipe_m2sPipe_payload_frameStart;
      controlStream_s2mPipe_m2sPipe_rData_rowEnd <= controlStream_s2mPipe_m2sPipe_payload_rowEnd;
      controlStream_s2mPipe_m2sPipe_rData_pipeValid <= controlStream_s2mPipe_m2sPipe_payload_pipeValid;
      controlStream_s2mPipe_m2sPipe_rData_firstRow <= controlStream_s2mPipe_m2sPipe_payload_firstRow;
      controlStream_s2mPipe_m2sPipe_rData_lastRow <= controlStream_s2mPipe_m2sPipe_payload_lastRow;
      controlStream_s2mPipe_m2sPipe_rData_finalResult <= controlStream_s2mPipe_m2sPipe_payload_finalResult;
      controlStream_s2mPipe_m2sPipe_rData_mainCompare <= controlStream_s2mPipe_m2sPipe_payload_mainCompare;
      controlStream_s2mPipe_m2sPipe_rData_counterCompare <= controlStream_s2mPipe_m2sPipe_payload_counterCompare;
      controlStream_s2mPipe_m2sPipe_rData_horizontalCompare <= controlStream_s2mPipe_m2sPipe_payload_horizontalCompare;
      controlStream_s2mPipe_m2sPipe_rData_verticalCompare <= controlStream_s2mPipe_m2sPipe_payload_verticalCompare;
      controlStream_s2mPipe_m2sPipe_rData_mainDiff <= controlStream_s2mPipe_m2sPipe_payload_mainDiff;
      controlStream_s2mPipe_m2sPipe_rData_counterDiff <= controlStream_s2mPipe_m2sPipe_payload_counterDiff;
      controlStream_s2mPipe_m2sPipe_rData_horizontalDiff <= controlStream_s2mPipe_m2sPipe_payload_horizontalDiff;
      controlStream_s2mPipe_m2sPipe_rData_verticalDiff <= controlStream_s2mPipe_m2sPipe_payload_verticalDiff;
      controlStream_s2mPipe_m2sPipe_rData_isHorizontalMin <= controlStream_s2mPipe_m2sPipe_payload_isHorizontalMin;
      controlStream_s2mPipe_m2sPipe_rData_minDiff <= controlStream_s2mPipe_m2sPipe_payload_minDiff;
      controlStream_s2mPipe_m2sPipe_rData_currentPosition <= controlStream_s2mPipe_m2sPipe_payload_currentPosition;
      controlStream_s2mPipe_m2sPipe_rData_nextPosition <= controlStream_s2mPipe_m2sPipe_payload_nextPosition;
      controlStream_s2mPipe_m2sPipe_rData_horizontalDirectionValid <= controlStream_s2mPipe_m2sPipe_payload_horizontalDirectionValid;
      controlStream_s2mPipe_m2sPipe_rData_verticalDirectionValid <= controlStream_s2mPipe_m2sPipe_payload_verticalDirectionValid;
      controlStream_s2mPipe_m2sPipe_rData_mainDirectionValid <= controlStream_s2mPipe_m2sPipe_payload_mainDirectionValid;
      controlStream_s2mPipe_m2sPipe_rData_counterDirectionValid <= controlStream_s2mPipe_m2sPipe_payload_counterDirectionValid;
      controlStream_s2mPipe_m2sPipe_rData_inValidMinDiff <= controlStream_s2mPipe_m2sPipe_payload_inValidMinDiff;
    end
    if(controlStream_s2mPipe_m2sPipe_m2sPipe_ready) begin
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_frameStart <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_frameStart;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_rowEnd <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_rowEnd;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_pipeValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_pipeValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_firstRow <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_firstRow;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_lastRow <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_lastRow;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_finalResult <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_finalResult;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_horizontalCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_horizontalCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_verticalCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_verticalCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_horizontalDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_horizontalDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_verticalDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_verticalDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_isHorizontalMin <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_isHorizontalMin;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_minDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_minDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_currentPosition <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_currentPosition;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_nextPosition <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_nextPosition;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_horizontalDirectionValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_horizontalDirectionValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_verticalDirectionValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_verticalDirectionValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainDirectionValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDirectionValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterDirectionValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDirectionValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_inValidMinDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_inValidMinDiff;
    end
    if(controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready) begin
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_frameStart <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_frameStart;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_rowEnd <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_rowEnd;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_pipeValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_pipeValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_firstRow <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_firstRow;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_lastRow <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_lastRow;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_finalResult <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_finalResult;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_horizontalCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_horizontalCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_verticalCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_verticalCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_horizontalDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_horizontalDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_verticalDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_verticalDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_isHorizontalMin <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_isHorizontalMin;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_minDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_minDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_currentPosition <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_currentPosition;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_nextPosition <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_nextPosition;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_horizontalDirectionValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_horizontalDirectionValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_verticalDirectionValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_verticalDirectionValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainDirectionValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainDirectionValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterDirectionValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterDirectionValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_inValidMinDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_inValidMinDiff;
    end
    if(readStage_mainOnePixelStream_ready) begin
      readStage_mainOnePixelStream_rData <= readStage_mainOnePixelStream_payload;
    end
    if(readStage_mainOnePixelStream_s2mPipe_ready) begin
      readStage_mainOnePixelStream_s2mPipe_rData <= readStage_mainOnePixelStream_s2mPipe_payload;
    end
    if(readStage_counterOnePixelStream_ready) begin
      readStage_counterOnePixelStream_rData <= readStage_counterOnePixelStream_payload;
    end
    if(readStage_counterOnePixelStream_s2mPipe_ready) begin
      readStage_counterOnePixelStream_s2mPipe_rData <= readStage_counterOnePixelStream_s2mPipe_payload;
    end
    if(readStage_mainTwoPixelStream_ready) begin
      readStage_mainTwoPixelStream_rData <= readStage_mainTwoPixelStream_payload;
    end
    if(readStage_mainTwoPixelStream_s2mPipe_ready) begin
      readStage_mainTwoPixelStream_s2mPipe_rData <= readStage_mainTwoPixelStream_s2mPipe_payload;
    end
    if(readStage_counterTwoPixelStream_ready) begin
      readStage_counterTwoPixelStream_rData <= readStage_counterTwoPixelStream_payload;
    end
    if(readStage_counterTwoPixelStream_s2mPipe_ready) begin
      readStage_counterTwoPixelStream_s2mPipe_rData <= readStage_counterTwoPixelStream_s2mPipe_payload;
    end
    if(readStage_mainThreePixelStream_ready) begin
      readStage_mainThreePixelStream_rData <= readStage_mainThreePixelStream_payload;
    end
    if(readStage_mainThreePixelStream_s2mPipe_ready) begin
      readStage_mainThreePixelStream_s2mPipe_rData <= readStage_mainThreePixelStream_s2mPipe_payload;
    end
    if(readStage_counterThreePixelStream_ready) begin
      readStage_counterThreePixelStream_rData <= readStage_counterThreePixelStream_payload;
    end
    if(readStage_counterThreePixelStream_s2mPipe_ready) begin
      readStage_counterThreePixelStream_s2mPipe_rData <= readStage_counterThreePixelStream_s2mPipe_payload;
    end
    if(readStage_mainOneValidStream_ready) begin
      readStage_mainOneValidStream_rData <= readStage_mainOneValidStream_payload;
    end
    if(readStage_mainOneValidStream_s2mPipe_ready) begin
      readStage_mainOneValidStream_s2mPipe_rData <= readStage_mainOneValidStream_s2mPipe_payload;
    end
    if(readStage_counterOneValidStream_ready) begin
      readStage_counterOneValidStream_rData <= readStage_counterOneValidStream_payload;
    end
    if(readStage_counterOneValidStream_s2mPipe_ready) begin
      readStage_counterOneValidStream_s2mPipe_rData <= readStage_counterOneValidStream_s2mPipe_payload;
    end
    if(readStage_mainTwoValidStream_ready) begin
      readStage_mainTwoValidStream_rData <= readStage_mainTwoValidStream_payload;
    end
    if(readStage_mainTwoValidStream_s2mPipe_ready) begin
      readStage_mainTwoValidStream_s2mPipe_rData <= readStage_mainTwoValidStream_s2mPipe_payload;
    end
    if(readStage_counterTwoValidStream_ready) begin
      readStage_counterTwoValidStream_rData <= readStage_counterTwoValidStream_payload;
    end
    if(readStage_counterTwoValidStream_s2mPipe_ready) begin
      readStage_counterTwoValidStream_s2mPipe_rData <= readStage_counterTwoValidStream_s2mPipe_payload;
    end
    if(readStage_mainThreeValidStream_ready) begin
      readStage_mainThreeValidStream_rData <= readStage_mainThreeValidStream_payload;
    end
    if(readStage_mainThreeValidStream_s2mPipe_ready) begin
      readStage_mainThreeValidStream_s2mPipe_rData <= readStage_mainThreeValidStream_s2mPipe_payload;
    end
    if(readStage_counterThreeValidStream_ready) begin
      readStage_counterThreeValidStream_rData <= readStage_counterThreeValidStream_payload;
    end
    if(readStage_counterThreeValidStream_s2mPipe_ready) begin
      readStage_counterThreeValidStream_s2mPipe_rData <= readStage_counterThreeValidStream_s2mPipe_payload;
    end
    if(readStage_controlPipe_translated_ready) begin
      readStage_controlPipe_translated_rData_frameStart <= readStage_controlPipe_translated_payload_frameStart;
      readStage_controlPipe_translated_rData_rowEnd <= readStage_controlPipe_translated_payload_rowEnd;
      readStage_controlPipe_translated_rData_pipeValid <= readStage_controlPipe_translated_payload_pipeValid;
      readStage_controlPipe_translated_rData_firstRow <= readStage_controlPipe_translated_payload_firstRow;
      readStage_controlPipe_translated_rData_lastRow <= readStage_controlPipe_translated_payload_lastRow;
      readStage_controlPipe_translated_rData_finalResult <= readStage_controlPipe_translated_payload_finalResult;
      readStage_controlPipe_translated_rData_mainCompare <= readStage_controlPipe_translated_payload_mainCompare;
      readStage_controlPipe_translated_rData_counterCompare <= readStage_controlPipe_translated_payload_counterCompare;
      readStage_controlPipe_translated_rData_horizontalCompare <= readStage_controlPipe_translated_payload_horizontalCompare;
      readStage_controlPipe_translated_rData_verticalCompare <= readStage_controlPipe_translated_payload_verticalCompare;
      readStage_controlPipe_translated_rData_mainDiff <= readStage_controlPipe_translated_payload_mainDiff;
      readStage_controlPipe_translated_rData_counterDiff <= readStage_controlPipe_translated_payload_counterDiff;
      readStage_controlPipe_translated_rData_horizontalDiff <= readStage_controlPipe_translated_payload_horizontalDiff;
      readStage_controlPipe_translated_rData_verticalDiff <= readStage_controlPipe_translated_payload_verticalDiff;
      readStage_controlPipe_translated_rData_isHorizontalMin <= readStage_controlPipe_translated_payload_isHorizontalMin;
      readStage_controlPipe_translated_rData_minDiff <= readStage_controlPipe_translated_payload_minDiff;
      readStage_controlPipe_translated_rData_currentPosition <= readStage_controlPipe_translated_payload_currentPosition;
      readStage_controlPipe_translated_rData_nextPosition <= readStage_controlPipe_translated_payload_nextPosition;
      readStage_controlPipe_translated_rData_horizontalDirectionValid <= readStage_controlPipe_translated_payload_horizontalDirectionValid;
      readStage_controlPipe_translated_rData_verticalDirectionValid <= readStage_controlPipe_translated_payload_verticalDirectionValid;
      readStage_controlPipe_translated_rData_mainDirectionValid <= readStage_controlPipe_translated_payload_mainDirectionValid;
      readStage_controlPipe_translated_rData_counterDirectionValid <= readStage_controlPipe_translated_payload_counterDirectionValid;
      readStage_controlPipe_translated_rData_inValidMinDiff <= readStage_controlPipe_translated_payload_inValidMinDiff;
    end
    if(readStage_controlPipe_translated_s2mPipe_ready) begin
      readStage_controlPipe_translated_s2mPipe_rData_frameStart <= readStage_controlPipe_translated_s2mPipe_payload_frameStart;
      readStage_controlPipe_translated_s2mPipe_rData_rowEnd <= readStage_controlPipe_translated_s2mPipe_payload_rowEnd;
      readStage_controlPipe_translated_s2mPipe_rData_pipeValid <= readStage_controlPipe_translated_s2mPipe_payload_pipeValid;
      readStage_controlPipe_translated_s2mPipe_rData_firstRow <= readStage_controlPipe_translated_s2mPipe_payload_firstRow;
      readStage_controlPipe_translated_s2mPipe_rData_lastRow <= readStage_controlPipe_translated_s2mPipe_payload_lastRow;
      readStage_controlPipe_translated_s2mPipe_rData_finalResult <= readStage_controlPipe_translated_s2mPipe_payload_finalResult;
      readStage_controlPipe_translated_s2mPipe_rData_mainCompare <= readStage_controlPipe_translated_s2mPipe_payload_mainCompare;
      readStage_controlPipe_translated_s2mPipe_rData_counterCompare <= readStage_controlPipe_translated_s2mPipe_payload_counterCompare;
      readStage_controlPipe_translated_s2mPipe_rData_horizontalCompare <= readStage_controlPipe_translated_s2mPipe_payload_horizontalCompare;
      readStage_controlPipe_translated_s2mPipe_rData_verticalCompare <= readStage_controlPipe_translated_s2mPipe_payload_verticalCompare;
      readStage_controlPipe_translated_s2mPipe_rData_mainDiff <= readStage_controlPipe_translated_s2mPipe_payload_mainDiff;
      readStage_controlPipe_translated_s2mPipe_rData_counterDiff <= readStage_controlPipe_translated_s2mPipe_payload_counterDiff;
      readStage_controlPipe_translated_s2mPipe_rData_horizontalDiff <= readStage_controlPipe_translated_s2mPipe_payload_horizontalDiff;
      readStage_controlPipe_translated_s2mPipe_rData_verticalDiff <= readStage_controlPipe_translated_s2mPipe_payload_verticalDiff;
      readStage_controlPipe_translated_s2mPipe_rData_isHorizontalMin <= readStage_controlPipe_translated_s2mPipe_payload_isHorizontalMin;
      readStage_controlPipe_translated_s2mPipe_rData_minDiff <= readStage_controlPipe_translated_s2mPipe_payload_minDiff;
      readStage_controlPipe_translated_s2mPipe_rData_currentPosition <= readStage_controlPipe_translated_s2mPipe_payload_currentPosition;
      readStage_controlPipe_translated_s2mPipe_rData_nextPosition <= readStage_controlPipe_translated_s2mPipe_payload_nextPosition;
      readStage_controlPipe_translated_s2mPipe_rData_horizontalDirectionValid <= readStage_controlPipe_translated_s2mPipe_payload_horizontalDirectionValid;
      readStage_controlPipe_translated_s2mPipe_rData_verticalDirectionValid <= readStage_controlPipe_translated_s2mPipe_payload_verticalDirectionValid;
      readStage_controlPipe_translated_s2mPipe_rData_mainDirectionValid <= readStage_controlPipe_translated_s2mPipe_payload_mainDirectionValid;
      readStage_controlPipe_translated_s2mPipe_rData_counterDirectionValid <= readStage_controlPipe_translated_s2mPipe_payload_counterDirectionValid;
      readStage_controlPipe_translated_s2mPipe_rData_inValidMinDiff <= readStage_controlPipe_translated_s2mPipe_payload_inValidMinDiff;
    end
    if(compareStage_mainOnePixelStream_ready) begin
      compareStage_mainOnePixelStream_rData <= compareStage_mainOnePixelStream_payload;
    end
    if(compareStage_mainOnePixelStream_s2mPipe_ready) begin
      compareStage_mainOnePixelStream_s2mPipe_rData <= compareStage_mainOnePixelStream_s2mPipe_payload;
    end
    if(compareStage_counterOnePixelStream_ready) begin
      compareStage_counterOnePixelStream_rData <= compareStage_counterOnePixelStream_payload;
    end
    if(compareStage_counterOnePixelStream_s2mPipe_ready) begin
      compareStage_counterOnePixelStream_s2mPipe_rData <= compareStage_counterOnePixelStream_s2mPipe_payload;
    end
    if(compareStage_mainTwoPixelStream_ready) begin
      compareStage_mainTwoPixelStream_rData <= compareStage_mainTwoPixelStream_payload;
    end
    if(compareStage_mainTwoPixelStream_s2mPipe_ready) begin
      compareStage_mainTwoPixelStream_s2mPipe_rData <= compareStage_mainTwoPixelStream_s2mPipe_payload;
    end
    if(compareStage_counterTwoPixelStream_ready) begin
      compareStage_counterTwoPixelStream_rData <= compareStage_counterTwoPixelStream_payload;
    end
    if(compareStage_counterTwoPixelStream_s2mPipe_ready) begin
      compareStage_counterTwoPixelStream_s2mPipe_rData <= compareStage_counterTwoPixelStream_s2mPipe_payload;
    end
    if(compareStage_mainThreePixelStream_ready) begin
      compareStage_mainThreePixelStream_rData <= compareStage_mainThreePixelStream_payload;
    end
    if(compareStage_mainThreePixelStream_s2mPipe_ready) begin
      compareStage_mainThreePixelStream_s2mPipe_rData <= compareStage_mainThreePixelStream_s2mPipe_payload;
    end
    if(compareStage_counterThreePixelStream_ready) begin
      compareStage_counterThreePixelStream_rData <= compareStage_counterThreePixelStream_payload;
    end
    if(compareStage_counterThreePixelStream_s2mPipe_ready) begin
      compareStage_counterThreePixelStream_s2mPipe_rData <= compareStage_counterThreePixelStream_s2mPipe_payload;
    end
    if(compareStage_mainOneValidStream_ready) begin
      compareStage_mainOneValidStream_rData <= compareStage_mainOneValidStream_payload;
    end
    if(compareStage_mainOneValidStream_s2mPipe_ready) begin
      compareStage_mainOneValidStream_s2mPipe_rData <= compareStage_mainOneValidStream_s2mPipe_payload;
    end
    if(compareStage_counterOneValidStream_ready) begin
      compareStage_counterOneValidStream_rData <= compareStage_counterOneValidStream_payload;
    end
    if(compareStage_counterOneValidStream_s2mPipe_ready) begin
      compareStage_counterOneValidStream_s2mPipe_rData <= compareStage_counterOneValidStream_s2mPipe_payload;
    end
    if(compareStage_mainTwoValidStream_ready) begin
      compareStage_mainTwoValidStream_rData <= compareStage_mainTwoValidStream_payload;
    end
    if(compareStage_mainTwoValidStream_s2mPipe_ready) begin
      compareStage_mainTwoValidStream_s2mPipe_rData <= compareStage_mainTwoValidStream_s2mPipe_payload;
    end
    if(compareStage_counterTwoValidStream_ready) begin
      compareStage_counterTwoValidStream_rData <= compareStage_counterTwoValidStream_payload;
    end
    if(compareStage_counterTwoValidStream_s2mPipe_ready) begin
      compareStage_counterTwoValidStream_s2mPipe_rData <= compareStage_counterTwoValidStream_s2mPipe_payload;
    end
    if(compareStage_mainThreeValidStream_ready) begin
      compareStage_mainThreeValidStream_rData <= compareStage_mainThreeValidStream_payload;
    end
    if(compareStage_mainThreeValidStream_s2mPipe_ready) begin
      compareStage_mainThreeValidStream_s2mPipe_rData <= compareStage_mainThreeValidStream_s2mPipe_payload;
    end
    if(compareStage_counterThreeValidStream_ready) begin
      compareStage_counterThreeValidStream_rData <= compareStage_counterThreeValidStream_payload;
    end
    if(compareStage_counterThreeValidStream_s2mPipe_ready) begin
      compareStage_counterThreeValidStream_s2mPipe_rData <= compareStage_counterThreeValidStream_s2mPipe_payload;
    end
    if(compareStage_controlPipe_translated_ready) begin
      compareStage_controlPipe_translated_rData_frameStart <= compareStage_controlPipe_translated_payload_frameStart;
      compareStage_controlPipe_translated_rData_rowEnd <= compareStage_controlPipe_translated_payload_rowEnd;
      compareStage_controlPipe_translated_rData_pipeValid <= compareStage_controlPipe_translated_payload_pipeValid;
      compareStage_controlPipe_translated_rData_firstRow <= compareStage_controlPipe_translated_payload_firstRow;
      compareStage_controlPipe_translated_rData_lastRow <= compareStage_controlPipe_translated_payload_lastRow;
      compareStage_controlPipe_translated_rData_finalResult <= compareStage_controlPipe_translated_payload_finalResult;
      compareStage_controlPipe_translated_rData_mainCompare <= compareStage_controlPipe_translated_payload_mainCompare;
      compareStage_controlPipe_translated_rData_counterCompare <= compareStage_controlPipe_translated_payload_counterCompare;
      compareStage_controlPipe_translated_rData_horizontalCompare <= compareStage_controlPipe_translated_payload_horizontalCompare;
      compareStage_controlPipe_translated_rData_verticalCompare <= compareStage_controlPipe_translated_payload_verticalCompare;
      compareStage_controlPipe_translated_rData_mainDiff <= compareStage_controlPipe_translated_payload_mainDiff;
      compareStage_controlPipe_translated_rData_counterDiff <= compareStage_controlPipe_translated_payload_counterDiff;
      compareStage_controlPipe_translated_rData_horizontalDiff <= compareStage_controlPipe_translated_payload_horizontalDiff;
      compareStage_controlPipe_translated_rData_verticalDiff <= compareStage_controlPipe_translated_payload_verticalDiff;
      compareStage_controlPipe_translated_rData_isHorizontalMin <= compareStage_controlPipe_translated_payload_isHorizontalMin;
      compareStage_controlPipe_translated_rData_minDiff <= compareStage_controlPipe_translated_payload_minDiff;
      compareStage_controlPipe_translated_rData_currentPosition <= compareStage_controlPipe_translated_payload_currentPosition;
      compareStage_controlPipe_translated_rData_nextPosition <= compareStage_controlPipe_translated_payload_nextPosition;
      compareStage_controlPipe_translated_rData_horizontalDirectionValid <= compareStage_controlPipe_translated_payload_horizontalDirectionValid;
      compareStage_controlPipe_translated_rData_verticalDirectionValid <= compareStage_controlPipe_translated_payload_verticalDirectionValid;
      compareStage_controlPipe_translated_rData_mainDirectionValid <= compareStage_controlPipe_translated_payload_mainDirectionValid;
      compareStage_controlPipe_translated_rData_counterDirectionValid <= compareStage_controlPipe_translated_payload_counterDirectionValid;
      compareStage_controlPipe_translated_rData_inValidMinDiff <= compareStage_controlPipe_translated_payload_inValidMinDiff;
    end
    if(compareStage_controlPipe_translated_s2mPipe_ready) begin
      compareStage_controlPipe_translated_s2mPipe_rData_frameStart <= compareStage_controlPipe_translated_s2mPipe_payload_frameStart;
      compareStage_controlPipe_translated_s2mPipe_rData_rowEnd <= compareStage_controlPipe_translated_s2mPipe_payload_rowEnd;
      compareStage_controlPipe_translated_s2mPipe_rData_pipeValid <= compareStage_controlPipe_translated_s2mPipe_payload_pipeValid;
      compareStage_controlPipe_translated_s2mPipe_rData_firstRow <= compareStage_controlPipe_translated_s2mPipe_payload_firstRow;
      compareStage_controlPipe_translated_s2mPipe_rData_lastRow <= compareStage_controlPipe_translated_s2mPipe_payload_lastRow;
      compareStage_controlPipe_translated_s2mPipe_rData_finalResult <= compareStage_controlPipe_translated_s2mPipe_payload_finalResult;
      compareStage_controlPipe_translated_s2mPipe_rData_mainCompare <= compareStage_controlPipe_translated_s2mPipe_payload_mainCompare;
      compareStage_controlPipe_translated_s2mPipe_rData_counterCompare <= compareStage_controlPipe_translated_s2mPipe_payload_counterCompare;
      compareStage_controlPipe_translated_s2mPipe_rData_horizontalCompare <= compareStage_controlPipe_translated_s2mPipe_payload_horizontalCompare;
      compareStage_controlPipe_translated_s2mPipe_rData_verticalCompare <= compareStage_controlPipe_translated_s2mPipe_payload_verticalCompare;
      compareStage_controlPipe_translated_s2mPipe_rData_mainDiff <= compareStage_controlPipe_translated_s2mPipe_payload_mainDiff;
      compareStage_controlPipe_translated_s2mPipe_rData_counterDiff <= compareStage_controlPipe_translated_s2mPipe_payload_counterDiff;
      compareStage_controlPipe_translated_s2mPipe_rData_horizontalDiff <= compareStage_controlPipe_translated_s2mPipe_payload_horizontalDiff;
      compareStage_controlPipe_translated_s2mPipe_rData_verticalDiff <= compareStage_controlPipe_translated_s2mPipe_payload_verticalDiff;
      compareStage_controlPipe_translated_s2mPipe_rData_isHorizontalMin <= compareStage_controlPipe_translated_s2mPipe_payload_isHorizontalMin;
      compareStage_controlPipe_translated_s2mPipe_rData_minDiff <= compareStage_controlPipe_translated_s2mPipe_payload_minDiff;
      compareStage_controlPipe_translated_s2mPipe_rData_currentPosition <= compareStage_controlPipe_translated_s2mPipe_payload_currentPosition;
      compareStage_controlPipe_translated_s2mPipe_rData_nextPosition <= compareStage_controlPipe_translated_s2mPipe_payload_nextPosition;
      compareStage_controlPipe_translated_s2mPipe_rData_horizontalDirectionValid <= compareStage_controlPipe_translated_s2mPipe_payload_horizontalDirectionValid;
      compareStage_controlPipe_translated_s2mPipe_rData_verticalDirectionValid <= compareStage_controlPipe_translated_s2mPipe_payload_verticalDirectionValid;
      compareStage_controlPipe_translated_s2mPipe_rData_mainDirectionValid <= compareStage_controlPipe_translated_s2mPipe_payload_mainDirectionValid;
      compareStage_controlPipe_translated_s2mPipe_rData_counterDirectionValid <= compareStage_controlPipe_translated_s2mPipe_payload_counterDirectionValid;
      compareStage_controlPipe_translated_s2mPipe_rData_inValidMinDiff <= compareStage_controlPipe_translated_s2mPipe_payload_inValidMinDiff;
    end
    if(diffStage_mainOnePixelStream_ready) begin
      diffStage_mainOnePixelStream_rData <= diffStage_mainOnePixelStream_payload;
    end
    if(diffStage_mainOnePixelStream_s2mPipe_ready) begin
      diffStage_mainOnePixelStream_s2mPipe_rData <= diffStage_mainOnePixelStream_s2mPipe_payload;
    end
    if(diffStage_counterOnePixelStream_ready) begin
      diffStage_counterOnePixelStream_rData <= diffStage_counterOnePixelStream_payload;
    end
    if(diffStage_counterOnePixelStream_s2mPipe_ready) begin
      diffStage_counterOnePixelStream_s2mPipe_rData <= diffStage_counterOnePixelStream_s2mPipe_payload;
    end
    if(diffStage_mainTwoPixelStream_ready) begin
      diffStage_mainTwoPixelStream_rData <= diffStage_mainTwoPixelStream_payload;
    end
    if(diffStage_mainTwoPixelStream_s2mPipe_ready) begin
      diffStage_mainTwoPixelStream_s2mPipe_rData <= diffStage_mainTwoPixelStream_s2mPipe_payload;
    end
    if(diffStage_counterTwoPixelStream_ready) begin
      diffStage_counterTwoPixelStream_rData <= diffStage_counterTwoPixelStream_payload;
    end
    if(diffStage_counterTwoPixelStream_s2mPipe_ready) begin
      diffStage_counterTwoPixelStream_s2mPipe_rData <= diffStage_counterTwoPixelStream_s2mPipe_payload;
    end
    if(diffStage_mainThreePixelStream_ready) begin
      diffStage_mainThreePixelStream_rData <= diffStage_mainThreePixelStream_payload;
    end
    if(diffStage_mainThreePixelStream_s2mPipe_ready) begin
      diffStage_mainThreePixelStream_s2mPipe_rData <= diffStage_mainThreePixelStream_s2mPipe_payload;
    end
    if(diffStage_counterThreePixelStream_ready) begin
      diffStage_counterThreePixelStream_rData <= diffStage_counterThreePixelStream_payload;
    end
    if(diffStage_counterThreePixelStream_s2mPipe_ready) begin
      diffStage_counterThreePixelStream_s2mPipe_rData <= diffStage_counterThreePixelStream_s2mPipe_payload;
    end
    if(diffStage_mainOneValidStream_ready) begin
      diffStage_mainOneValidStream_rData <= diffStage_mainOneValidStream_payload;
    end
    if(diffStage_mainOneValidStream_s2mPipe_ready) begin
      diffStage_mainOneValidStream_s2mPipe_rData <= diffStage_mainOneValidStream_s2mPipe_payload;
    end
    if(diffStage_counterOneValidStream_ready) begin
      diffStage_counterOneValidStream_rData <= diffStage_counterOneValidStream_payload;
    end
    if(diffStage_counterOneValidStream_s2mPipe_ready) begin
      diffStage_counterOneValidStream_s2mPipe_rData <= diffStage_counterOneValidStream_s2mPipe_payload;
    end
    if(diffStage_mainTwoValidStream_ready) begin
      diffStage_mainTwoValidStream_rData <= diffStage_mainTwoValidStream_payload;
    end
    if(diffStage_mainTwoValidStream_s2mPipe_ready) begin
      diffStage_mainTwoValidStream_s2mPipe_rData <= diffStage_mainTwoValidStream_s2mPipe_payload;
    end
    if(diffStage_counterTwoValidStream_ready) begin
      diffStage_counterTwoValidStream_rData <= diffStage_counterTwoValidStream_payload;
    end
    if(diffStage_counterTwoValidStream_s2mPipe_ready) begin
      diffStage_counterTwoValidStream_s2mPipe_rData <= diffStage_counterTwoValidStream_s2mPipe_payload;
    end
    if(diffStage_mainThreeValidStream_ready) begin
      diffStage_mainThreeValidStream_rData <= diffStage_mainThreeValidStream_payload;
    end
    if(diffStage_mainThreeValidStream_s2mPipe_ready) begin
      diffStage_mainThreeValidStream_s2mPipe_rData <= diffStage_mainThreeValidStream_s2mPipe_payload;
    end
    if(diffStage_counterThreeValidStream_ready) begin
      diffStage_counterThreeValidStream_rData <= diffStage_counterThreeValidStream_payload;
    end
    if(diffStage_counterThreeValidStream_s2mPipe_ready) begin
      diffStage_counterThreeValidStream_s2mPipe_rData <= diffStage_counterThreeValidStream_s2mPipe_payload;
    end
    if(resultStage_controlPipeBeforePipe_ready) begin
      resultStage_controlPipeBeforePipe_rData_frameStart <= resultStage_controlPipeBeforePipe_payload_frameStart;
      resultStage_controlPipeBeforePipe_rData_rowEnd <= resultStage_controlPipeBeforePipe_payload_rowEnd;
      resultStage_controlPipeBeforePipe_rData_pipeValid <= resultStage_controlPipeBeforePipe_payload_pipeValid;
      resultStage_controlPipeBeforePipe_rData_firstRow <= resultStage_controlPipeBeforePipe_payload_firstRow;
      resultStage_controlPipeBeforePipe_rData_lastRow <= resultStage_controlPipeBeforePipe_payload_lastRow;
      resultStage_controlPipeBeforePipe_rData_finalResult <= resultStage_controlPipeBeforePipe_payload_finalResult;
      resultStage_controlPipeBeforePipe_rData_mainCompare <= resultStage_controlPipeBeforePipe_payload_mainCompare;
      resultStage_controlPipeBeforePipe_rData_counterCompare <= resultStage_controlPipeBeforePipe_payload_counterCompare;
      resultStage_controlPipeBeforePipe_rData_horizontalCompare <= resultStage_controlPipeBeforePipe_payload_horizontalCompare;
      resultStage_controlPipeBeforePipe_rData_verticalCompare <= resultStage_controlPipeBeforePipe_payload_verticalCompare;
      resultStage_controlPipeBeforePipe_rData_mainDiff <= resultStage_controlPipeBeforePipe_payload_mainDiff;
      resultStage_controlPipeBeforePipe_rData_counterDiff <= resultStage_controlPipeBeforePipe_payload_counterDiff;
      resultStage_controlPipeBeforePipe_rData_horizontalDiff <= resultStage_controlPipeBeforePipe_payload_horizontalDiff;
      resultStage_controlPipeBeforePipe_rData_verticalDiff <= resultStage_controlPipeBeforePipe_payload_verticalDiff;
      resultStage_controlPipeBeforePipe_rData_isHorizontalMin <= resultStage_controlPipeBeforePipe_payload_isHorizontalMin;
      resultStage_controlPipeBeforePipe_rData_minDiff <= resultStage_controlPipeBeforePipe_payload_minDiff;
      resultStage_controlPipeBeforePipe_rData_currentPosition <= resultStage_controlPipeBeforePipe_payload_currentPosition;
      resultStage_controlPipeBeforePipe_rData_nextPosition <= resultStage_controlPipeBeforePipe_payload_nextPosition;
      resultStage_controlPipeBeforePipe_rData_horizontalDirectionValid <= resultStage_controlPipeBeforePipe_payload_horizontalDirectionValid;
      resultStage_controlPipeBeforePipe_rData_verticalDirectionValid <= resultStage_controlPipeBeforePipe_payload_verticalDirectionValid;
      resultStage_controlPipeBeforePipe_rData_mainDirectionValid <= resultStage_controlPipeBeforePipe_payload_mainDirectionValid;
      resultStage_controlPipeBeforePipe_rData_counterDirectionValid <= resultStage_controlPipeBeforePipe_payload_counterDirectionValid;
      resultStage_controlPipeBeforePipe_rData_inValidMinDiff <= resultStage_controlPipeBeforePipe_payload_inValidMinDiff;
    end
    if(resultStage_controlPipeBeforePipe_s2mPipe_ready) begin
      resultStage_controlPipeBeforePipe_s2mPipe_rData_frameStart <= resultStage_controlPipeBeforePipe_s2mPipe_payload_frameStart;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_rowEnd <= resultStage_controlPipeBeforePipe_s2mPipe_payload_rowEnd;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_pipeValid <= resultStage_controlPipeBeforePipe_s2mPipe_payload_pipeValid;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_firstRow <= resultStage_controlPipeBeforePipe_s2mPipe_payload_firstRow;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_lastRow <= resultStage_controlPipeBeforePipe_s2mPipe_payload_lastRow;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_finalResult <= resultStage_controlPipeBeforePipe_s2mPipe_payload_finalResult;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_mainCompare <= resultStage_controlPipeBeforePipe_s2mPipe_payload_mainCompare;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_counterCompare <= resultStage_controlPipeBeforePipe_s2mPipe_payload_counterCompare;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_horizontalCompare <= resultStage_controlPipeBeforePipe_s2mPipe_payload_horizontalCompare;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_verticalCompare <= resultStage_controlPipeBeforePipe_s2mPipe_payload_verticalCompare;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_mainDiff <= resultStage_controlPipeBeforePipe_s2mPipe_payload_mainDiff;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_counterDiff <= resultStage_controlPipeBeforePipe_s2mPipe_payload_counterDiff;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_horizontalDiff <= resultStage_controlPipeBeforePipe_s2mPipe_payload_horizontalDiff;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_verticalDiff <= resultStage_controlPipeBeforePipe_s2mPipe_payload_verticalDiff;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_isHorizontalMin <= resultStage_controlPipeBeforePipe_s2mPipe_payload_isHorizontalMin;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_minDiff <= resultStage_controlPipeBeforePipe_s2mPipe_payload_minDiff;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_currentPosition <= resultStage_controlPipeBeforePipe_s2mPipe_payload_currentPosition;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_nextPosition <= resultStage_controlPipeBeforePipe_s2mPipe_payload_nextPosition;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_horizontalDirectionValid <= resultStage_controlPipeBeforePipe_s2mPipe_payload_horizontalDirectionValid;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_verticalDirectionValid <= resultStage_controlPipeBeforePipe_s2mPipe_payload_verticalDirectionValid;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_mainDirectionValid <= resultStage_controlPipeBeforePipe_s2mPipe_payload_mainDirectionValid;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_counterDirectionValid <= resultStage_controlPipeBeforePipe_s2mPipe_payload_counterDirectionValid;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_inValidMinDiff <= resultStage_controlPipeBeforePipe_s2mPipe_payload_inValidMinDiff;
    end
    if(resultStage_pixelStream_ready) begin
      resultStage_pixelStream_rData <= resultStage_pixelStream_payload;
    end
    if(resultStage_pixelStream_s2mPipe_ready) begin
      resultStage_pixelStream_s2mPipe_rData <= resultStage_pixelStream_s2mPipe_payload;
    end
    if(pixelsStream_ready) begin
      pixelsStream_rData_pixel <= pixelsStream_payload_pixel;
      pixelsStream_rData_frameStart <= pixelsStream_payload_frameStart;
      pixelsStream_rData_rowEnd <= pixelsStream_payload_rowEnd;
    end
    if(pixelsStream_s2mPipe_ready) begin
      pixelsStream_s2mPipe_rData_pixel <= pixelsStream_s2mPipe_payload_pixel;
      pixelsStream_s2mPipe_rData_frameStart <= pixelsStream_s2mPipe_payload_frameStart;
      pixelsStream_s2mPipe_rData_rowEnd <= pixelsStream_s2mPipe_payload_rowEnd;
    end
  end


endmodule

module SuperResolutionPart2_1 (
  input               pixelsIn_valid,
  output reg          pixelsIn_ready,
  input      [7:0]    pixelsIn_payload_pixel,
  input               pixelsIn_payload_frameStart,
  input               pixelsIn_payload_rowEnd,
  input               startIn,
  input               inpThreeDoneIn,
  output reg          pixelsOut_valid,
  input               pixelsOut_ready,
  output reg [7:0]    pixelsOut_payload_pixel,
  output reg          pixelsOut_payload_frameStart,
  output reg          pixelsOut_payload_rowEnd,
  output reg          pixelsOut_payload_inpValid,
  output reg          startOut,
  output reg          inpTwoDoneOut,
  input      [7:0]    thresholdIn,
  input      [9:0]    widthIn,
  input      [9:0]    heightIn,
  input               clk,
  input               resetn
);
  localparam controlStateMachine_enumDef_4_BOOT = 3'd0;
  localparam controlStateMachine_enumDef_4_HOLD = 3'd1;
  localparam controlStateMachine_enumDef_4_PASS = 3'd2;
  localparam controlStateMachine_enumDef_4_ONCE = 3'd3;
  localparam controlStateMachine_enumDef_4_TWICE = 3'd4;

  reg        [7:0]    CICC1851_lineBufferOne_port1;
  reg        [7:0]    CICC1851_lineBufferOne_port2;
  reg        [7:0]    CICC1851_lineBufferTwo_port1;
  reg        [7:0]    CICC1851_lineBufferTwo_port2;
  reg        [7:0]    CICC1851_lineBufferOdd_port1;
  wire                diffStage_controlPipe_fork_io_input_ready;
  wire                diffStage_controlPipe_fork_io_outputs_0_valid;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_frameStart;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_rowEnd;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_passMode;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_passValid;
  wire       [2:0]    diffStage_controlPipe_fork_io_outputs_0_payload_onceMode;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_onceValid;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_mainCompare;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_counterCompare;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_payload_mainDiff;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_payload_counterDiff;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_twiceCompValid;
  wire       [2:0]    diffStage_controlPipe_fork_io_outputs_0_payload_twiceMode;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_inpValidFlag;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_oddValid;
  wire                diffStage_controlPipe_fork_io_outputs_1_valid;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_frameStart;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_rowEnd;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_passMode;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_passValid;
  wire       [2:0]    diffStage_controlPipe_fork_io_outputs_1_payload_onceMode;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_onceValid;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_mainCompare;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_counterCompare;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_twiceCompValid;
  wire       [2:0]    diffStage_controlPipe_fork_io_outputs_1_payload_twiceMode;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_inpValidFlag;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_oddValid;
  wire       [10:0]   CICC1851_bufferRowCount_valueNext;
  wire       [0:0]    CICC1851_bufferRowCount_valueNext_1;
  wire       [10:0]   CICC1851_bufferWAddr_valueNext;
  wire       [0:0]    CICC1851_bufferWAddr_valueNext_1;
  wire       [11:0]   CICC1851_outPixelAddr_valueNext;
  wire       [0:0]    CICC1851_outPixelAddr_valueNext_1;
  wire       [11:0]   CICC1851_outRowCount_valueNext;
  wire       [0:0]    CICC1851_outRowCount_valueNext_1;
  wire       [11:0]   CICC1851_alreadySendRow_valueNext;
  wire       [0:0]    CICC1851_alreadySendRow_valueNext_1;
  wire       [11:0]   CICC1851_alreadySendCountInRow_valueNext;
  wire       [0:0]    CICC1851_alreadySendCountInRow_valueNext_1;
  wire       [11:0]   CICC1851_mainAddrOne;
  wire       [11:0]   CICC1851_counterAddrOne;
  wire       [11:0]   CICC1851_mainAddrTwo;
  wire       [11:0]   CICC1851_counterAddrTwo;
  wire       [11:0]   CICC1851_oddAddr;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l181;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l181_1;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l181_2;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l182;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l182_1;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l182_2;
  wire       [10:0]   CICC1851_when_SuperResolutionPart2_l195;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l218;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l234;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l234_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l234_2;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l235;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l235_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l235_2;
  wire       [7:0]    CICC1851_lineBufferOne_port;
  wire                CICC1851_lineBufferOne_port_1;
  wire       [7:0]    CICC1851_lineBufferOdd_port;
  wire                CICC1851_lineBufferOdd_port_1;
  wire       [7:0]    CICC1851_lineBufferTwo_port;
  wire                CICC1851_lineBufferTwo_port_1;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_1;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_2;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_3;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_4;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_5;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_6;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_7;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_8;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_9;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_10;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_11;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_12;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_13;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_14;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_15;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_16;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_17;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_18;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_19;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l763;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l763_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l763_2;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l764;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l764_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l764_2;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l783;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l785;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l787;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l789;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l793;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l796;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l799;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l802;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l560;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l560_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l602;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l602_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l602_2;
  wire       [2:0]    CICC1851_when_SuperResolutionPart2_l602_3;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l603;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l603_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l605;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l605_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l605_2;
  wire       [2:0]    CICC1851_when_SuperResolutionPart2_l605_3;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l606;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l606_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l606_2;
  wire       [1:0]    CICC1851_when_SuperResolutionPart2_l606_3;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l609;
  wire       [11:0]   CICC1851_mainAddrOne_1;
  wire       [11:0]   CICC1851_mainAddrOne_2;
  wire       [11:0]   CICC1851_mainAddrTwo_1;
  wire       [11:0]   CICC1851_mainAddrTwo_2;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l667;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l667_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l667_2;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l667_3;
  wire       [1:0]    CICC1851_when_SuperResolutionPart2_l667_4;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l668;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l668_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l668_2;
  wire       [1:0]    CICC1851_when_SuperResolutionPart2_l668_3;
  wire       [11:0]   CICC1851_mainAddrOne_3;
  wire       [11:0]   CICC1851_mainAddrOne_4;
  wire       [11:0]   CICC1851_mainAddrTwo_3;
  wire       [11:0]   CICC1851_mainAddrTwo_4;
  wire       [1:0]    CICC1851_controls_onceMode;
  wire       [1:0]    CICC1851_controls_onceMode_1;
  wire       [11:0]   CICC1851_mainAddrOne_5;
  wire       [11:0]   CICC1851_mainAddrOne_6;
  wire       [11:0]   CICC1851_counterAddrOne_1;
  wire       [11:0]   CICC1851_counterAddrOne_2;
  wire       [11:0]   CICC1851_counterAddrOne_3;
  wire       [11:0]   CICC1851_counterAddrOne_4;
  wire       [0:0]    CICC1851_controls_onceMode_2;
  wire       [11:0]   CICC1851_mainAddrTwo_5;
  wire       [11:0]   CICC1851_mainAddrTwo_6;
  wire       [11:0]   CICC1851_counterAddrTwo_1;
  wire       [11:0]   CICC1851_counterAddrTwo_2;
  wire       [11:0]   CICC1851_counterAddrTwo_3;
  wire       [11:0]   CICC1851_counterAddrTwo_4;
  wire       [11:0]   CICC1851_mainAddrOne_7;
  wire       [11:0]   CICC1851_mainAddrOne_8;
  wire       [11:0]   CICC1851_mainAddrOne_9;
  wire       [11:0]   CICC1851_mainAddrOne_10;
  wire       [12:0]   CICC1851_counterAddrOne_5;
  wire       [12:0]   CICC1851_counterAddrOne_6;
  wire       [12:0]   CICC1851_counterAddrOne_7;
  wire       [1:0]    CICC1851_counterAddrOne_8;
  wire       [1:0]    CICC1851_controls_twiceMode;
  wire       [11:0]   CICC1851_mainAddrTwo_7;
  wire       [11:0]   CICC1851_mainAddrTwo_8;
  wire       [1:0]    CICC1851_controls_twiceMode_1;
  wire       [11:0]   CICC1851_mainAddrTwo_9;
  wire       [11:0]   CICC1851_mainAddrTwo_10;
  wire       [12:0]   CICC1851_counterAddrTwo_5;
  wire       [12:0]   CICC1851_counterAddrTwo_6;
  wire       [12:0]   CICC1851_counterAddrTwo_7;
  wire       [1:0]    CICC1851_counterAddrTwo_8;
  wire       [11:0]   CICC1851_mainAddrOne_11;
  wire       [11:0]   CICC1851_mainAddrOne_12;
  wire       [11:0]   CICC1851_counterAddrTwo_9;
  wire       [11:0]   CICC1851_counterAddrTwo_10;
  wire       [11:0]   CICC1851_mainAddrTwo_11;
  wire       [11:0]   CICC1851_mainAddrTwo_12;
  wire       [11:0]   CICC1851_counterAddrOne_9;
  wire       [11:0]   CICC1851_counterAddrOne_10;
  wire       [12:0]   CICC1851_mainAddrTwo_13;
  wire       [12:0]   CICC1851_mainAddrTwo_14;
  wire       [12:0]   CICC1851_mainAddrTwo_15;
  wire       [1:0]    CICC1851_mainAddrTwo_16;
  wire       [12:0]   CICC1851_counterAddrOne_11;
  wire       [12:0]   CICC1851_counterAddrOne_12;
  wire       [12:0]   CICC1851_counterAddrOne_13;
  wire       [1:0]    CICC1851_counterAddrOne_14;
  wire       [0:0]    CICC1851_controls_twiceMode_2;
  wire       [11:0]   CICC1851_mainAddrTwo_17;
  wire       [11:0]   CICC1851_mainAddrTwo_18;
  wire       [11:0]   CICC1851_counterAddrOne_15;
  wire       [11:0]   CICC1851_counterAddrOne_16;
  wire       [11:0]   CICC1851_mainAddrOne_13;
  wire       [11:0]   CICC1851_mainAddrOne_14;
  wire       [11:0]   CICC1851_counterAddrTwo_11;
  wire       [11:0]   CICC1851_counterAddrTwo_12;
  wire       [12:0]   CICC1851_mainAddrOne_15;
  wire       [12:0]   CICC1851_mainAddrOne_16;
  wire       [12:0]   CICC1851_mainAddrOne_17;
  wire       [1:0]    CICC1851_mainAddrOne_18;
  wire       [12:0]   CICC1851_counterAddrTwo_13;
  wire       [12:0]   CICC1851_counterAddrTwo_14;
  wire       [12:0]   CICC1851_counterAddrTwo_15;
  wire       [1:0]    CICC1851_counterAddrTwo_16;
  reg                 inpTwoDone;
  reg                 startIn_regNext;
  wire                when_SuperResolutionPart2_l40;
  reg                 readDone;
  wire                when_SuperResolutionPart2_l43;
  reg                 startRead;
  wire                when_SuperResolutionPart2_l46;
  wire                when_SuperResolutionPart2_l46_1;
  reg                 slaveStart;
  wire                pixelsIn_fire;
  wire                when_SuperResolutionPart2_l49;
  wire                when_SuperResolutionPart2_l49_1;
  reg                 frameStart;
  reg        [7:0]    inpThreshold;
  reg        [9:0]    bmpWidth;
  reg        [9:0]    bmpHeight;
  reg                 holdBuffer;
  wire                when_SuperResolutionPart2_l64;
  reg                 writeDone;
  wire                when_SuperResolutionPart2_l67;
  reg                 bufferRowCount_willIncrement;
  reg                 bufferRowCount_willClear;
  reg        [10:0]   bufferRowCount_valueNext;
  reg        [10:0]   bufferRowCount_value;
  wire                bufferRowCount_willOverflowIfInc;
  wire                bufferRowCount_willOverflow;
  reg                 bufferReuse;
  reg                 bufferEnable;
  wire                when_SuperResolutionPart2_l76;
  wire                when_SuperResolutionPart2_l76_1;
  reg        [1:0]    bufferSwitch;
  reg                 nextRowBuffer;
  wire                when_SuperResolutionPart2_l82;
  reg                 bufferWAddr_willIncrement;
  reg                 bufferWAddr_willClear;
  reg        [10:0]   bufferWAddr_valueNext;
  reg        [10:0]   bufferWAddr_value;
  wire                bufferWAddr_willOverflowIfInc;
  wire                bufferWAddr_willOverflow;
  reg                 outPixelAddr_willIncrement;
  reg                 outPixelAddr_willClear;
  reg        [11:0]   outPixelAddr_valueNext;
  reg        [11:0]   outPixelAddr_value;
  wire                outPixelAddr_willOverflowIfInc;
  wire                outPixelAddr_willOverflow;
  reg                 outRowCount_willIncrement;
  reg                 outRowCount_willClear;
  reg        [11:0]   outRowCount_valueNext;
  reg        [11:0]   outRowCount_value;
  wire                outRowCount_willOverflowIfInc;
  wire                outRowCount_willOverflow;
  reg                 alreadySendRow_willIncrement;
  reg                 alreadySendRow_willClear;
  reg        [11:0]   alreadySendRow_valueNext;
  reg        [11:0]   alreadySendRow_value;
  wire                alreadySendRow_willOverflowIfInc;
  wire                alreadySendRow_willOverflow;
  reg                 alreadySendCountInRow_willIncrement;
  reg                 alreadySendCountInRow_willClear;
  reg        [11:0]   alreadySendCountInRow_valueNext;
  reg        [11:0]   alreadySendCountInRow_value;
  wire                alreadySendCountInRow_willOverflowIfInc;
  wire                alreadySendCountInRow_willOverflow;
  reg                 alreadyReachRowEnd;
  reg                 alreadyReachFinalRow;
  reg                 outReachRowEnd;
  reg                 outReachFinalRow;
  reg                 bufferReachRowEnd;
  reg                 bufferReachFinalRow;
  reg                 oddBufferRow;
  reg                 startIn_regNext_1;
  wire                when_SuperResolutionPart2_l106;
  reg                 zeroInFourOutPixelAddr;
  reg                 startIn_regNext_2;
  wire                when_SuperResolutionPart2_l108;
  reg                 oneInFourOutPixelAddr;
  reg                 startIn_regNext_3;
  wire                when_SuperResolutionPart2_l109;
  reg                 twoInFourOutPixelAddr;
  reg                 startIn_regNext_4;
  wire                when_SuperResolutionPart2_l110;
  reg                 threeInFourOutPixelAddr;
  reg                 startIn_regNext_5;
  wire                when_SuperResolutionPart2_l111;
  reg                 zeroInFourOutRow;
  reg                 startIn_regNext_6;
  wire                when_SuperResolutionPart2_l113;
  reg                 oneInFourOutRow;
  reg                 startIn_regNext_7;
  wire                when_SuperResolutionPart2_l114;
  reg                 twoInFourOutRow;
  reg                 startIn_regNext_8;
  wire                when_SuperResolutionPart2_l115;
  reg                 threeInFourOutRow;
  reg                 startIn_regNext_9;
  wire                when_SuperResolutionPart2_l116;
  wire       [2:0]    currentState;
  reg                 willHoldToTwice;
  reg                 startIn_regNext_10;
  wire                when_SuperResolutionPart2_l120;
  reg                 willPassToHoldCaseOne;
  reg                 startIn_regNext_11;
  wire                when_SuperResolutionPart2_l121;
  reg                 willPassToHoldCaseTwo;
  reg                 startIn_regNext_12;
  wire                when_SuperResolutionPart2_l122;
  reg                 holdWillPassToHoldCaseTwo;
  reg                 startIn_regNext_13;
  wire                when_SuperResolutionPart2_l123;
  reg                 willOnceToHoldCaseOne;
  reg                 startIn_regNext_14;
  wire                when_SuperResolutionPart2_l124;
  reg                 willOnceToHoldCaseTwo;
  reg                 startIn_regNext_15;
  wire                when_SuperResolutionPart2_l125;
  reg                 willOnceToHoldCaseThree;
  reg                 startIn_regNext_16;
  wire                when_SuperResolutionPart2_l126;
  wire                when_SuperResolutionPart2_l134;
  reg        [10:0]   mainAddrOne;
  reg        [10:0]   counterAddrOne;
  reg        [10:0]   mainAddrTwo;
  reg        [10:0]   counterAddrTwo;
  wire       [10:0]   oddAddr;
  wire                validStream_valid;
  reg                 validStream_ready;
  wire                controlStream_valid;
  wire                controlStream_ready;
  wire                controlStream_payload_frameStart;
  wire                controlStream_payload_rowEnd;
  wire                controlStream_payload_passMode;
  wire                controlStream_payload_passValid;
  wire       [2:0]    controlStream_payload_onceMode;
  wire                controlStream_payload_onceValid;
  wire                controlStream_payload_mainCompare;
  wire                controlStream_payload_counterCompare;
  wire       [7:0]    controlStream_payload_mainDiff;
  wire       [7:0]    controlStream_payload_counterDiff;
  wire                controlStream_payload_twiceCompValid;
  wire       [2:0]    controlStream_payload_twiceMode;
  wire                controlStream_payload_inpValidFlag;
  wire                controlStream_payload_oddValid;
  reg                 controls_frameStart;
  reg                 controls_rowEnd;
  reg                 controls_passMode;
  reg                 controls_passValid;
  reg        [2:0]    controls_onceMode;
  reg                 controls_onceValid;
  wire                controls_mainCompare;
  wire                controls_counterCompare;
  wire       [7:0]    controls_mainDiff;
  wire       [7:0]    controls_counterDiff;
  reg                 controls_twiceCompValid;
  reg        [2:0]    controls_twiceMode;
  reg                 controls_inpValidFlag;
  reg                 controls_oddValid;
  wire       [31:0]   CICC1851_controls_frameStart;
  wire                mainAddrOneStream_valid;
  wire                mainAddrOneStream_ready;
  wire       [10:0]   mainAddrOneStream_payload;
  wire                counterAddrOneStream_valid;
  wire                counterAddrOneStream_ready;
  wire       [10:0]   counterAddrOneStream_payload;
  wire                mainAddrTwoStream_valid;
  wire                mainAddrTwoStream_ready;
  wire       [10:0]   mainAddrTwoStream_payload;
  wire                counterAddrTwoStream_valid;
  wire                counterAddrTwoStream_ready;
  wire       [10:0]   counterAddrTwoStream_payload;
  wire                oddAddrStream_valid;
  wire                oddAddrStream_ready;
  wire       [10:0]   oddAddrStream_payload;
  wire                pixelsIn_s2mPipe_valid;
  reg                 pixelsIn_s2mPipe_ready;
  wire       [7:0]    pixelsIn_s2mPipe_payload_pixel;
  wire                pixelsIn_s2mPipe_payload_frameStart;
  wire                pixelsIn_s2mPipe_payload_rowEnd;
  reg                 pixelsIn_rValid;
  reg        [7:0]    pixelsIn_rData_pixel;
  reg                 pixelsIn_rData_frameStart;
  reg                 pixelsIn_rData_rowEnd;
  wire                pixelsIn_s2mPipe_m2sPipe_valid;
  wire                pixelsIn_s2mPipe_m2sPipe_ready;
  wire       [7:0]    pixelsIn_s2mPipe_m2sPipe_payload_pixel;
  wire                pixelsIn_s2mPipe_m2sPipe_payload_frameStart;
  wire                pixelsIn_s2mPipe_m2sPipe_payload_rowEnd;
  reg                 pixelsIn_s2mPipe_rValid;
  reg        [7:0]    pixelsIn_s2mPipe_rData_pixel;
  reg                 pixelsIn_s2mPipe_rData_frameStart;
  reg                 pixelsIn_s2mPipe_rData_rowEnd;
  wire                when_Stream_l368;
  wire                passPixels_valid;
  wire                passPixels_ready;
  wire       [7:0]    passPixels_payload_pixel;
  wire                passPixels_payload_frameStart;
  wire                passPixels_payload_rowEnd;
  wire                passPixels_fire;
  wire                when_SuperResolutionPart2_l181;
  wire                passPixels_fire_1;
  wire                when_SuperResolutionPart2_l182;
  wire                passPixels_fire_2;
  wire                when_SuperResolutionPart2_l185;
  wire                when_SuperResolutionPart2_l195;
  wire                passPixels_fire_3;
  wire                when_SuperResolutionPart2_l200;
  wire                when_SuperResolutionPart2_l201;
  wire                passPixels_fire_4;
  wire                when_SuperResolutionPart2_l207;
  wire                when_SuperResolutionPart2_l208;
  wire                when_SuperResolutionPart2_l212;
  wire                controlStream_fire;
  wire                when_SuperResolutionPart2_l218;
  wire                when_SuperResolutionPart2_l220;
  wire                passPixels_fire_5;
  wire                when_SuperResolutionPart2_l224;
  wire                pixelsOut_fire;
  wire                when_SuperResolutionPart2_l234;
  wire                pixelsOut_fire_1;
  wire                when_SuperResolutionPart2_l235;
  wire                pixelsOut_fire_2;
  wire                pixelsOut_fire_3;
  wire                when_SuperResolutionPart2_l246;
  wire                passPixels_fire_6;
  wire                passPixels_fire_7;
  wire                passPixels_fire_8;
  wire                passPixels_fire_9;
  wire                passPixels_fire_10;
  wire                controlStream_fire_1;
  wire                pushing;
  wire                passPixels_fire_11;
  wire                controlStream_fire_2;
  wire                poping;
  wire                passPixels_fire_12;
  wire                controlStream_fire_3;
  wire                pushAndPoping;
  wire                mainAddrOneStream_s2mPipe_valid;
  reg                 mainAddrOneStream_s2mPipe_ready;
  wire       [10:0]   mainAddrOneStream_s2mPipe_payload;
  reg                 mainAddrOneStream_rValid;
  reg        [10:0]   mainAddrOneStream_rData;
  wire                mainAddrOneStream_s2mPipe_m2sPipe_valid;
  wire                mainAddrOneStream_s2mPipe_m2sPipe_ready;
  wire       [10:0]   mainAddrOneStream_s2mPipe_m2sPipe_payload;
  reg                 mainAddrOneStream_s2mPipe_rValid;
  reg        [10:0]   mainAddrOneStream_s2mPipe_rData;
  wire                when_Stream_l368_1;
  wire                CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_mainOnePixelStream_payload;
  reg                 CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_1;
  reg                 CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_mainOnePixelStream_payload_1;
  wire                readStage_mainOnePixelStream_valid;
  wire                readStage_mainOnePixelStream_ready;
  wire       [7:0]    readStage_mainOnePixelStream_payload;
  reg                 CICC1851_readStage_mainOnePixelStream_valid;
  reg        [7:0]    CICC1851_readStage_mainOnePixelStream_payload_2;
  wire                when_Stream_l368_2;
  wire                counterAddrOneStream_s2mPipe_valid;
  reg                 counterAddrOneStream_s2mPipe_ready;
  wire       [10:0]   counterAddrOneStream_s2mPipe_payload;
  reg                 counterAddrOneStream_rValid;
  reg        [10:0]   counterAddrOneStream_rData;
  wire                counterAddrOneStream_s2mPipe_m2sPipe_valid;
  wire                counterAddrOneStream_s2mPipe_m2sPipe_ready;
  wire       [10:0]   counterAddrOneStream_s2mPipe_m2sPipe_payload;
  reg                 counterAddrOneStream_s2mPipe_rValid;
  reg        [10:0]   counterAddrOneStream_s2mPipe_rData;
  wire                when_Stream_l368_3;
  wire                CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_counterOnePixelStream_payload;
  reg                 CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_2;
  reg                 CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_counterOnePixelStream_payload_1;
  wire                readStage_counterOnePixelStream_valid;
  wire                readStage_counterOnePixelStream_ready;
  wire       [7:0]    readStage_counterOnePixelStream_payload;
  reg                 CICC1851_readStage_counterOnePixelStream_valid;
  reg        [7:0]    CICC1851_readStage_counterOnePixelStream_payload_2;
  wire                when_Stream_l368_4;
  wire                mainAddrTwoStream_s2mPipe_valid;
  reg                 mainAddrTwoStream_s2mPipe_ready;
  wire       [10:0]   mainAddrTwoStream_s2mPipe_payload;
  reg                 mainAddrTwoStream_rValid;
  reg        [10:0]   mainAddrTwoStream_rData;
  wire                mainAddrTwoStream_s2mPipe_m2sPipe_valid;
  wire                mainAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire       [10:0]   mainAddrTwoStream_s2mPipe_m2sPipe_payload;
  reg                 mainAddrTwoStream_s2mPipe_rValid;
  reg        [10:0]   mainAddrTwoStream_s2mPipe_rData;
  wire                when_Stream_l368_5;
  wire                CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_mainTwoPixelStream_payload;
  reg                 CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_3;
  reg                 CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_mainTwoPixelStream_payload_1;
  wire                readStage_mainTwoPixelStream_valid;
  wire                readStage_mainTwoPixelStream_ready;
  wire       [7:0]    readStage_mainTwoPixelStream_payload;
  reg                 CICC1851_readStage_mainTwoPixelStream_valid;
  reg        [7:0]    CICC1851_readStage_mainTwoPixelStream_payload_2;
  wire                when_Stream_l368_6;
  wire                counterAddrTwoStream_s2mPipe_valid;
  reg                 counterAddrTwoStream_s2mPipe_ready;
  wire       [10:0]   counterAddrTwoStream_s2mPipe_payload;
  reg                 counterAddrTwoStream_rValid;
  reg        [10:0]   counterAddrTwoStream_rData;
  wire                counterAddrTwoStream_s2mPipe_m2sPipe_valid;
  wire                counterAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire       [10:0]   counterAddrTwoStream_s2mPipe_m2sPipe_payload;
  reg                 counterAddrTwoStream_s2mPipe_rValid;
  reg        [10:0]   counterAddrTwoStream_s2mPipe_rData;
  wire                when_Stream_l368_7;
  wire                CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_counterTwoPixelStream_payload;
  reg                 CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_4;
  reg                 CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_counterTwoPixelStream_payload_1;
  wire                readStage_counterTwoPixelStream_valid;
  wire                readStage_counterTwoPixelStream_ready;
  wire       [7:0]    readStage_counterTwoPixelStream_payload;
  reg                 CICC1851_readStage_counterTwoPixelStream_valid;
  reg        [7:0]    CICC1851_readStage_counterTwoPixelStream_payload_2;
  wire                when_Stream_l368_8;
  wire                oddAddrStream_s2mPipe_valid;
  reg                 oddAddrStream_s2mPipe_ready;
  wire       [10:0]   oddAddrStream_s2mPipe_payload;
  reg                 oddAddrStream_rValid;
  reg        [10:0]   oddAddrStream_rData;
  wire                oddAddrStream_s2mPipe_m2sPipe_valid;
  wire                oddAddrStream_s2mPipe_m2sPipe_ready;
  wire       [10:0]   oddAddrStream_s2mPipe_m2sPipe_payload;
  reg                 oddAddrStream_s2mPipe_rValid;
  reg        [10:0]   oddAddrStream_s2mPipe_rData;
  wire                when_Stream_l368_9;
  wire                CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_oddRowPixelStream_payload;
  reg                 CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_5;
  reg                 CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_oddRowPixelStream_payload_1;
  wire                readStage_oddRowPixelStream_valid;
  wire                readStage_oddRowPixelStream_ready;
  wire       [7:0]    readStage_oddRowPixelStream_payload;
  reg                 CICC1851_readStage_oddRowPixelStream_valid;
  reg        [7:0]    CICC1851_readStage_oddRowPixelStream_payload_2;
  wire                when_Stream_l368_10;
  wire                controlStream_s2mPipe_valid;
  reg                 controlStream_s2mPipe_ready;
  wire                controlStream_s2mPipe_payload_frameStart;
  wire                controlStream_s2mPipe_payload_rowEnd;
  wire                controlStream_s2mPipe_payload_passMode;
  wire                controlStream_s2mPipe_payload_passValid;
  wire       [2:0]    controlStream_s2mPipe_payload_onceMode;
  wire                controlStream_s2mPipe_payload_onceValid;
  wire                controlStream_s2mPipe_payload_mainCompare;
  wire                controlStream_s2mPipe_payload_counterCompare;
  wire       [7:0]    controlStream_s2mPipe_payload_mainDiff;
  wire       [7:0]    controlStream_s2mPipe_payload_counterDiff;
  wire                controlStream_s2mPipe_payload_twiceCompValid;
  wire       [2:0]    controlStream_s2mPipe_payload_twiceMode;
  wire                controlStream_s2mPipe_payload_inpValidFlag;
  wire                controlStream_s2mPipe_payload_oddValid;
  reg                 controlStream_rValid;
  reg                 controlStream_rData_frameStart;
  reg                 controlStream_rData_rowEnd;
  reg                 controlStream_rData_passMode;
  reg                 controlStream_rData_passValid;
  reg        [2:0]    controlStream_rData_onceMode;
  reg                 controlStream_rData_onceValid;
  reg                 controlStream_rData_mainCompare;
  reg                 controlStream_rData_counterCompare;
  reg        [7:0]    controlStream_rData_mainDiff;
  reg        [7:0]    controlStream_rData_counterDiff;
  reg                 controlStream_rData_twiceCompValid;
  reg        [2:0]    controlStream_rData_twiceMode;
  reg                 controlStream_rData_inpValidFlag;
  reg                 controlStream_rData_oddValid;
  wire                controlStream_s2mPipe_m2sPipe_valid;
  reg                 controlStream_s2mPipe_m2sPipe_ready;
  wire                controlStream_s2mPipe_m2sPipe_payload_frameStart;
  wire                controlStream_s2mPipe_m2sPipe_payload_rowEnd;
  wire                controlStream_s2mPipe_m2sPipe_payload_passMode;
  wire                controlStream_s2mPipe_m2sPipe_payload_passValid;
  wire       [2:0]    controlStream_s2mPipe_m2sPipe_payload_onceMode;
  wire                controlStream_s2mPipe_m2sPipe_payload_onceValid;
  wire                controlStream_s2mPipe_m2sPipe_payload_mainCompare;
  wire                controlStream_s2mPipe_m2sPipe_payload_counterCompare;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_payload_mainDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_payload_counterDiff;
  wire                controlStream_s2mPipe_m2sPipe_payload_twiceCompValid;
  wire       [2:0]    controlStream_s2mPipe_m2sPipe_payload_twiceMode;
  wire                controlStream_s2mPipe_m2sPipe_payload_inpValidFlag;
  wire                controlStream_s2mPipe_m2sPipe_payload_oddValid;
  reg                 controlStream_s2mPipe_rValid;
  reg                 controlStream_s2mPipe_rData_frameStart;
  reg                 controlStream_s2mPipe_rData_rowEnd;
  reg                 controlStream_s2mPipe_rData_passMode;
  reg                 controlStream_s2mPipe_rData_passValid;
  reg        [2:0]    controlStream_s2mPipe_rData_onceMode;
  reg                 controlStream_s2mPipe_rData_onceValid;
  reg                 controlStream_s2mPipe_rData_mainCompare;
  reg                 controlStream_s2mPipe_rData_counterCompare;
  reg        [7:0]    controlStream_s2mPipe_rData_mainDiff;
  reg        [7:0]    controlStream_s2mPipe_rData_counterDiff;
  reg                 controlStream_s2mPipe_rData_twiceCompValid;
  reg        [2:0]    controlStream_s2mPipe_rData_twiceMode;
  reg                 controlStream_s2mPipe_rData_inpValidFlag;
  reg                 controlStream_s2mPipe_rData_oddValid;
  wire                when_Stream_l368_11;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_valid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_ready;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_frameStart;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_rowEnd;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passMode;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passValid;
  wire       [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceMode;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceValid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainCompare;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterCompare;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDiff;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceCompValid;
  wire       [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceMode;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_inpValidFlag;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_oddValid;
  reg                 controlStream_s2mPipe_m2sPipe_rValid;
  reg                 controlStream_s2mPipe_m2sPipe_rData_frameStart;
  reg                 controlStream_s2mPipe_m2sPipe_rData_rowEnd;
  reg                 controlStream_s2mPipe_m2sPipe_rData_passMode;
  reg                 controlStream_s2mPipe_m2sPipe_rData_passValid;
  reg        [2:0]    controlStream_s2mPipe_m2sPipe_rData_onceMode;
  reg                 controlStream_s2mPipe_m2sPipe_rData_onceValid;
  reg                 controlStream_s2mPipe_m2sPipe_rData_mainCompare;
  reg                 controlStream_s2mPipe_m2sPipe_rData_counterCompare;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_rData_mainDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_rData_counterDiff;
  reg                 controlStream_s2mPipe_m2sPipe_rData_twiceCompValid;
  reg        [2:0]    controlStream_s2mPipe_m2sPipe_rData_twiceMode;
  reg                 controlStream_s2mPipe_m2sPipe_rData_inpValidFlag;
  reg                 controlStream_s2mPipe_m2sPipe_rData_oddValid;
  wire                when_Stream_l368_12;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_valid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_frameStart;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_rowEnd;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_passMode;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_passValid;
  wire       [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_onceMode;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_onceValid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainCompare;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterCompare;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterDiff;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_twiceCompValid;
  wire       [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_twiceMode;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_inpValidFlag;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_oddValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_frameStart;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_rowEnd;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_passMode;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_passValid;
  reg        [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_onceMode;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_onceValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainCompare;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterCompare;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterDiff;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_twiceCompValid;
  reg        [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_twiceMode;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_inpValidFlag;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_oddValid;
  wire                readStage_controlPipe_valid;
  wire                readStage_controlPipe_ready;
  wire                readStage_controlPipe_payload_frameStart;
  wire                readStage_controlPipe_payload_rowEnd;
  wire                readStage_controlPipe_payload_passMode;
  wire                readStage_controlPipe_payload_passValid;
  wire       [2:0]    readStage_controlPipe_payload_onceMode;
  wire                readStage_controlPipe_payload_onceValid;
  wire                readStage_controlPipe_payload_mainCompare;
  wire                readStage_controlPipe_payload_counterCompare;
  wire       [7:0]    readStage_controlPipe_payload_mainDiff;
  wire       [7:0]    readStage_controlPipe_payload_counterDiff;
  wire                readStage_controlPipe_payload_twiceCompValid;
  wire       [2:0]    readStage_controlPipe_payload_twiceMode;
  wire                readStage_controlPipe_payload_inpValidFlag;
  wire                readStage_controlPipe_payload_oddValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_frameStart;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_rowEnd;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_passMode;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_passValid;
  reg        [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_onceMode;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_onceValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainCompare;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterCompare;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterDiff;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_twiceCompValid;
  reg        [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_twiceMode;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_inpValidFlag;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_oddValid;
  wire                when_Stream_l368_13;
  wire                readStage_mainOnePixelStream_s2mPipe_valid;
  reg                 readStage_mainOnePixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_mainOnePixelStream_s2mPipe_payload;
  reg                 readStage_mainOnePixelStream_rValid;
  reg        [7:0]    readStage_mainOnePixelStream_rData;
  wire                compareStage_mainOnePixelStream_valid;
  wire                compareStage_mainOnePixelStream_ready;
  wire       [7:0]    compareStage_mainOnePixelStream_payload;
  reg                 readStage_mainOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_mainOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_14;
  wire                readStage_counterOnePixelStream_s2mPipe_valid;
  reg                 readStage_counterOnePixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_counterOnePixelStream_s2mPipe_payload;
  reg                 readStage_counterOnePixelStream_rValid;
  reg        [7:0]    readStage_counterOnePixelStream_rData;
  wire                compareStage_counterOnePixelStream_valid;
  wire                compareStage_counterOnePixelStream_ready;
  wire       [7:0]    compareStage_counterOnePixelStream_payload;
  reg                 readStage_counterOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_counterOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_15;
  wire                readStage_mainTwoPixelStream_s2mPipe_valid;
  reg                 readStage_mainTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_mainTwoPixelStream_s2mPipe_payload;
  reg                 readStage_mainTwoPixelStream_rValid;
  reg        [7:0]    readStage_mainTwoPixelStream_rData;
  wire                compareStage_mainTwoPixelStream_valid;
  wire                compareStage_mainTwoPixelStream_ready;
  wire       [7:0]    compareStage_mainTwoPixelStream_payload;
  reg                 readStage_mainTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_mainTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_16;
  wire                readStage_counterTwoPixelStream_s2mPipe_valid;
  reg                 readStage_counterTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_counterTwoPixelStream_s2mPipe_payload;
  reg                 readStage_counterTwoPixelStream_rValid;
  reg        [7:0]    readStage_counterTwoPixelStream_rData;
  wire                compareStage_counterTwoPixelStream_valid;
  wire                compareStage_counterTwoPixelStream_ready;
  wire       [7:0]    compareStage_counterTwoPixelStream_payload;
  reg                 readStage_counterTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_counterTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_17;
  wire                readStage_oddRowPixelStream_s2mPipe_valid;
  reg                 readStage_oddRowPixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_oddRowPixelStream_s2mPipe_payload;
  reg                 readStage_oddRowPixelStream_rValid;
  reg        [7:0]    readStage_oddRowPixelStream_rData;
  wire                compareStage_oddRowPixelStream_valid;
  wire                compareStage_oddRowPixelStream_ready;
  wire       [7:0]    compareStage_oddRowPixelStream_payload;
  reg                 readStage_oddRowPixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_oddRowPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_18;
  reg                 CICC1851_readStage_controlPipe_translated_payload_mainCompare;
  reg                 CICC1851_readStage_controlPipe_translated_payload_counterCompare;
  wire                when_SuperResolutionPart2_l290;
  wire                when_SuperResolutionPart2_l294;
  wire                when_SuperResolutionPart2_l298;
  wire                when_SuperResolutionPart2_l302;
  wire                when_SuperResolutionPart2_l313;
  wire                when_SuperResolutionPart2_l315;
  wire                when_SuperResolutionPart2_l319;
  wire                when_SuperResolutionPart2_l321;
  wire                when_SuperResolutionPart2_l326;
  wire                when_SuperResolutionPart2_l331;
  wire                readStage_controlPipe_translated_valid;
  wire                readStage_controlPipe_translated_ready;
  wire                readStage_controlPipe_translated_payload_frameStart;
  wire                readStage_controlPipe_translated_payload_rowEnd;
  wire                readStage_controlPipe_translated_payload_passMode;
  wire                readStage_controlPipe_translated_payload_passValid;
  wire       [2:0]    readStage_controlPipe_translated_payload_onceMode;
  wire                readStage_controlPipe_translated_payload_onceValid;
  wire                readStage_controlPipe_translated_payload_mainCompare;
  wire                readStage_controlPipe_translated_payload_counterCompare;
  wire       [7:0]    readStage_controlPipe_translated_payload_mainDiff;
  wire       [7:0]    readStage_controlPipe_translated_payload_counterDiff;
  wire                readStage_controlPipe_translated_payload_twiceCompValid;
  wire       [2:0]    readStage_controlPipe_translated_payload_twiceMode;
  wire                readStage_controlPipe_translated_payload_inpValidFlag;
  wire                readStage_controlPipe_translated_payload_oddValid;
  wire                readStage_controlPipe_translated_s2mPipe_valid;
  reg                 readStage_controlPipe_translated_s2mPipe_ready;
  wire                readStage_controlPipe_translated_s2mPipe_payload_frameStart;
  wire                readStage_controlPipe_translated_s2mPipe_payload_rowEnd;
  wire                readStage_controlPipe_translated_s2mPipe_payload_passMode;
  wire                readStage_controlPipe_translated_s2mPipe_payload_passValid;
  wire       [2:0]    readStage_controlPipe_translated_s2mPipe_payload_onceMode;
  wire                readStage_controlPipe_translated_s2mPipe_payload_onceValid;
  wire                readStage_controlPipe_translated_s2mPipe_payload_mainCompare;
  wire                readStage_controlPipe_translated_s2mPipe_payload_counterCompare;
  wire       [7:0]    readStage_controlPipe_translated_s2mPipe_payload_mainDiff;
  wire       [7:0]    readStage_controlPipe_translated_s2mPipe_payload_counterDiff;
  wire                readStage_controlPipe_translated_s2mPipe_payload_twiceCompValid;
  wire       [2:0]    readStage_controlPipe_translated_s2mPipe_payload_twiceMode;
  wire                readStage_controlPipe_translated_s2mPipe_payload_inpValidFlag;
  wire                readStage_controlPipe_translated_s2mPipe_payload_oddValid;
  reg                 readStage_controlPipe_translated_rValid;
  reg                 readStage_controlPipe_translated_rData_frameStart;
  reg                 readStage_controlPipe_translated_rData_rowEnd;
  reg                 readStage_controlPipe_translated_rData_passMode;
  reg                 readStage_controlPipe_translated_rData_passValid;
  reg        [2:0]    readStage_controlPipe_translated_rData_onceMode;
  reg                 readStage_controlPipe_translated_rData_onceValid;
  reg                 readStage_controlPipe_translated_rData_mainCompare;
  reg                 readStage_controlPipe_translated_rData_counterCompare;
  reg        [7:0]    readStage_controlPipe_translated_rData_mainDiff;
  reg        [7:0]    readStage_controlPipe_translated_rData_counterDiff;
  reg                 readStage_controlPipe_translated_rData_twiceCompValid;
  reg        [2:0]    readStage_controlPipe_translated_rData_twiceMode;
  reg                 readStage_controlPipe_translated_rData_inpValidFlag;
  reg                 readStage_controlPipe_translated_rData_oddValid;
  wire                compareStage_controlPipe_valid;
  wire                compareStage_controlPipe_ready;
  wire                compareStage_controlPipe_payload_frameStart;
  wire                compareStage_controlPipe_payload_rowEnd;
  wire                compareStage_controlPipe_payload_passMode;
  wire                compareStage_controlPipe_payload_passValid;
  wire       [2:0]    compareStage_controlPipe_payload_onceMode;
  wire                compareStage_controlPipe_payload_onceValid;
  wire                compareStage_controlPipe_payload_mainCompare;
  wire                compareStage_controlPipe_payload_counterCompare;
  wire       [7:0]    compareStage_controlPipe_payload_mainDiff;
  wire       [7:0]    compareStage_controlPipe_payload_counterDiff;
  wire                compareStage_controlPipe_payload_twiceCompValid;
  wire       [2:0]    compareStage_controlPipe_payload_twiceMode;
  wire                compareStage_controlPipe_payload_inpValidFlag;
  wire                compareStage_controlPipe_payload_oddValid;
  reg                 readStage_controlPipe_translated_s2mPipe_rValid;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_frameStart;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_rowEnd;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_passMode;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_passValid;
  reg        [2:0]    readStage_controlPipe_translated_s2mPipe_rData_onceMode;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_onceValid;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_mainCompare;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_counterCompare;
  reg        [7:0]    readStage_controlPipe_translated_s2mPipe_rData_mainDiff;
  reg        [7:0]    readStage_controlPipe_translated_s2mPipe_rData_counterDiff;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_twiceCompValid;
  reg        [2:0]    readStage_controlPipe_translated_s2mPipe_rData_twiceMode;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_inpValidFlag;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_oddValid;
  wire                when_Stream_l368_19;
  wire                compareStage_mainOnePixelStream_s2mPipe_valid;
  reg                 compareStage_mainOnePixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_mainOnePixelStream_s2mPipe_payload;
  reg                 compareStage_mainOnePixelStream_rValid;
  reg        [7:0]    compareStage_mainOnePixelStream_rData;
  wire                diffStage_mainOnePixelStream_valid;
  wire                diffStage_mainOnePixelStream_ready;
  wire       [7:0]    diffStage_mainOnePixelStream_payload;
  reg                 compareStage_mainOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_mainOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_20;
  wire                compareStage_counterOnePixelStream_s2mPipe_valid;
  reg                 compareStage_counterOnePixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_counterOnePixelStream_s2mPipe_payload;
  reg                 compareStage_counterOnePixelStream_rValid;
  reg        [7:0]    compareStage_counterOnePixelStream_rData;
  wire                diffStage_counterOnePixelStream_valid;
  wire                diffStage_counterOnePixelStream_ready;
  wire       [7:0]    diffStage_counterOnePixelStream_payload;
  reg                 compareStage_counterOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_counterOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_21;
  wire                compareStage_mainTwoPixelStream_s2mPipe_valid;
  reg                 compareStage_mainTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_mainTwoPixelStream_s2mPipe_payload;
  reg                 compareStage_mainTwoPixelStream_rValid;
  reg        [7:0]    compareStage_mainTwoPixelStream_rData;
  wire                diffStage_mainTwoPixelStream_valid;
  wire                diffStage_mainTwoPixelStream_ready;
  wire       [7:0]    diffStage_mainTwoPixelStream_payload;
  reg                 compareStage_mainTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_mainTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_22;
  wire                compareStage_counterTwoPixelStream_s2mPipe_valid;
  reg                 compareStage_counterTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_counterTwoPixelStream_s2mPipe_payload;
  reg                 compareStage_counterTwoPixelStream_rValid;
  reg        [7:0]    compareStage_counterTwoPixelStream_rData;
  wire                diffStage_counterTwoPixelStream_valid;
  wire                diffStage_counterTwoPixelStream_ready;
  wire       [7:0]    diffStage_counterTwoPixelStream_payload;
  reg                 compareStage_counterTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_counterTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_23;
  wire                compareStage_oddRowPixelStream_s2mPipe_valid;
  reg                 compareStage_oddRowPixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_oddRowPixelStream_s2mPipe_payload;
  reg                 compareStage_oddRowPixelStream_rValid;
  reg        [7:0]    compareStage_oddRowPixelStream_rData;
  wire                diffStage_oddRowPixelStream_valid;
  wire                diffStage_oddRowPixelStream_ready;
  wire       [7:0]    diffStage_oddRowPixelStream_payload;
  reg                 compareStage_oddRowPixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_oddRowPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_24;
  reg        [7:0]    CICC1851_compareStage_controlPipe_translated_payload_mainDiff;
  reg        [7:0]    CICC1851_compareStage_controlPipe_translated_payload_counterDiff;
  wire                compareStage_controlPipe_translated_valid;
  wire                compareStage_controlPipe_translated_ready;
  wire                compareStage_controlPipe_translated_payload_frameStart;
  wire                compareStage_controlPipe_translated_payload_rowEnd;
  wire                compareStage_controlPipe_translated_payload_passMode;
  wire                compareStage_controlPipe_translated_payload_passValid;
  wire       [2:0]    compareStage_controlPipe_translated_payload_onceMode;
  wire                compareStage_controlPipe_translated_payload_onceValid;
  wire                compareStage_controlPipe_translated_payload_mainCompare;
  wire                compareStage_controlPipe_translated_payload_counterCompare;
  wire       [7:0]    compareStage_controlPipe_translated_payload_mainDiff;
  wire       [7:0]    compareStage_controlPipe_translated_payload_counterDiff;
  wire                compareStage_controlPipe_translated_payload_twiceCompValid;
  wire       [2:0]    compareStage_controlPipe_translated_payload_twiceMode;
  wire                compareStage_controlPipe_translated_payload_inpValidFlag;
  wire                compareStage_controlPipe_translated_payload_oddValid;
  wire                compareStage_controlPipe_translated_s2mPipe_valid;
  reg                 compareStage_controlPipe_translated_s2mPipe_ready;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_frameStart;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_rowEnd;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_passMode;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_passValid;
  wire       [2:0]    compareStage_controlPipe_translated_s2mPipe_payload_onceMode;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_onceValid;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_mainCompare;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_counterCompare;
  wire       [7:0]    compareStage_controlPipe_translated_s2mPipe_payload_mainDiff;
  wire       [7:0]    compareStage_controlPipe_translated_s2mPipe_payload_counterDiff;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_twiceCompValid;
  wire       [2:0]    compareStage_controlPipe_translated_s2mPipe_payload_twiceMode;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_inpValidFlag;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_oddValid;
  reg                 compareStage_controlPipe_translated_rValid;
  reg                 compareStage_controlPipe_translated_rData_frameStart;
  reg                 compareStage_controlPipe_translated_rData_rowEnd;
  reg                 compareStage_controlPipe_translated_rData_passMode;
  reg                 compareStage_controlPipe_translated_rData_passValid;
  reg        [2:0]    compareStage_controlPipe_translated_rData_onceMode;
  reg                 compareStage_controlPipe_translated_rData_onceValid;
  reg                 compareStage_controlPipe_translated_rData_mainCompare;
  reg                 compareStage_controlPipe_translated_rData_counterCompare;
  reg        [7:0]    compareStage_controlPipe_translated_rData_mainDiff;
  reg        [7:0]    compareStage_controlPipe_translated_rData_counterDiff;
  reg                 compareStage_controlPipe_translated_rData_twiceCompValid;
  reg        [2:0]    compareStage_controlPipe_translated_rData_twiceMode;
  reg                 compareStage_controlPipe_translated_rData_inpValidFlag;
  reg                 compareStage_controlPipe_translated_rData_oddValid;
  wire                diffStage_controlPipe_valid;
  wire                diffStage_controlPipe_ready;
  wire                diffStage_controlPipe_payload_frameStart;
  wire                diffStage_controlPipe_payload_rowEnd;
  wire                diffStage_controlPipe_payload_passMode;
  wire                diffStage_controlPipe_payload_passValid;
  wire       [2:0]    diffStage_controlPipe_payload_onceMode;
  wire                diffStage_controlPipe_payload_onceValid;
  wire                diffStage_controlPipe_payload_mainCompare;
  wire                diffStage_controlPipe_payload_counterCompare;
  wire       [7:0]    diffStage_controlPipe_payload_mainDiff;
  wire       [7:0]    diffStage_controlPipe_payload_counterDiff;
  wire                diffStage_controlPipe_payload_twiceCompValid;
  wire       [2:0]    diffStage_controlPipe_payload_twiceMode;
  wire                diffStage_controlPipe_payload_inpValidFlag;
  wire                diffStage_controlPipe_payload_oddValid;
  reg                 compareStage_controlPipe_translated_s2mPipe_rValid;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_frameStart;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_rowEnd;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_passMode;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_passValid;
  reg        [2:0]    compareStage_controlPipe_translated_s2mPipe_rData_onceMode;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_onceValid;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_mainCompare;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_counterCompare;
  reg        [7:0]    compareStage_controlPipe_translated_s2mPipe_rData_mainDiff;
  reg        [7:0]    compareStage_controlPipe_translated_s2mPipe_rData_counterDiff;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_twiceCompValid;
  reg        [2:0]    compareStage_controlPipe_translated_s2mPipe_rData_twiceMode;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_inpValidFlag;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_oddValid;
  wire                when_Stream_l368_25;
  wire                diffStage_mainOnePixelStream_s2mPipe_valid;
  reg                 diffStage_mainOnePixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_mainOnePixelStream_s2mPipe_payload;
  reg                 diffStage_mainOnePixelStream_rValid;
  reg        [7:0]    diffStage_mainOnePixelStream_rData;
  wire                resultStage_mainOnePixelStream_valid;
  wire                resultStage_mainOnePixelStream_ready;
  wire       [7:0]    resultStage_mainOnePixelStream_payload;
  reg                 diffStage_mainOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_mainOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_26;
  wire                diffStage_counterOnePixelStream_s2mPipe_valid;
  reg                 diffStage_counterOnePixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_counterOnePixelStream_s2mPipe_payload;
  reg                 diffStage_counterOnePixelStream_rValid;
  reg        [7:0]    diffStage_counterOnePixelStream_rData;
  wire                resultStage_counterOnePixelStream_valid;
  wire                resultStage_counterOnePixelStream_ready;
  wire       [7:0]    resultStage_counterOnePixelStream_payload;
  reg                 diffStage_counterOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_counterOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_27;
  wire                diffStage_mainTwoPixelStream_s2mPipe_valid;
  reg                 diffStage_mainTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_mainTwoPixelStream_s2mPipe_payload;
  reg                 diffStage_mainTwoPixelStream_rValid;
  reg        [7:0]    diffStage_mainTwoPixelStream_rData;
  wire                resultStage_mainTwoPixelStream_valid;
  wire                resultStage_mainTwoPixelStream_ready;
  wire       [7:0]    resultStage_mainTwoPixelStream_payload;
  reg                 diffStage_mainTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_mainTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_28;
  wire                diffStage_counterTwoPixelStream_s2mPipe_valid;
  reg                 diffStage_counterTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_counterTwoPixelStream_s2mPipe_payload;
  reg                 diffStage_counterTwoPixelStream_rValid;
  reg        [7:0]    diffStage_counterTwoPixelStream_rData;
  wire                resultStage_counterTwoPixelStream_valid;
  wire                resultStage_counterTwoPixelStream_ready;
  wire       [7:0]    resultStage_counterTwoPixelStream_payload;
  reg                 diffStage_counterTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_counterTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_29;
  wire                diffStage_oddRowPixelStream_s2mPipe_valid;
  reg                 diffStage_oddRowPixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_oddRowPixelStream_s2mPipe_payload;
  reg                 diffStage_oddRowPixelStream_rValid;
  reg        [7:0]    diffStage_oddRowPixelStream_rData;
  wire                resultStage_oddRowPixelStream_valid;
  wire                resultStage_oddRowPixelStream_ready;
  wire       [7:0]    resultStage_oddRowPixelStream_payload;
  reg                 diffStage_oddRowPixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_oddRowPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_30;
  wire       [2:0]    CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceMode;
  wire                CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceValid;
  wire       [7:0]    CICC1851_when_SuperResolutionPart2_l419;
  wire       [7:0]    CICC1851_when_SuperResolutionPart2_l428;
  wire                CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceCompValid;
  wire       [2:0]    CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceMode;
  reg                 CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag;
  wire                when_SuperResolutionPart2_l419;
  wire                when_SuperResolutionPart2_l420;
  wire                when_SuperResolutionPart2_l421;
  wire                when_SuperResolutionPart2_l422;
  wire                when_SuperResolutionPart2_l428;
  wire                when_SuperResolutionPart2_l429;
  wire                when_SuperResolutionPart2_l430;
  wire                when_SuperResolutionPart2_l431;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_valid;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_ready;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_payload_frameStart;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_payload_rowEnd;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_payload_passMode;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_payload_passValid;
  wire       [2:0]    diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceMode;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceValid;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_payload_mainCompare;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_payload_counterCompare;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_translated_payload_mainDiff;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_translated_payload_counterDiff;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceCompValid;
  wire       [2:0]    diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceMode;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_payload_oddValid;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_valid;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_ready;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_frameStart;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_rowEnd;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_passMode;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_passValid;
  wire       [2:0]    diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_onceMode;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_onceValid;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_mainCompare;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_counterCompare;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_mainDiff;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_counterDiff;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_twiceCompValid;
  wire       [2:0]    diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_twiceMode;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_inpValidFlag;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_oddValid;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_rValid;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_rData_frameStart;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_rData_rowEnd;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_rData_passMode;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_rData_passValid;
  reg        [2:0]    diffStage_controlPipe_fork_io_outputs_0_translated_rData_onceMode;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_rData_onceValid;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_rData_mainCompare;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_rData_counterCompare;
  reg        [7:0]    diffStage_controlPipe_fork_io_outputs_0_translated_rData_mainDiff;
  reg        [7:0]    diffStage_controlPipe_fork_io_outputs_0_translated_rData_counterDiff;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_rData_twiceCompValid;
  reg        [2:0]    diffStage_controlPipe_fork_io_outputs_0_translated_rData_twiceMode;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_rData_inpValidFlag;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_rData_oddValid;
  wire                resultStage_controlPipe_valid;
  wire                resultStage_controlPipe_ready;
  wire                resultStage_controlPipe_payload_frameStart;
  wire                resultStage_controlPipe_payload_rowEnd;
  wire                resultStage_controlPipe_payload_passMode;
  wire                resultStage_controlPipe_payload_passValid;
  wire       [2:0]    resultStage_controlPipe_payload_onceMode;
  wire                resultStage_controlPipe_payload_onceValid;
  wire                resultStage_controlPipe_payload_mainCompare;
  wire                resultStage_controlPipe_payload_counterCompare;
  wire       [7:0]    resultStage_controlPipe_payload_mainDiff;
  wire       [7:0]    resultStage_controlPipe_payload_counterDiff;
  wire                resultStage_controlPipe_payload_twiceCompValid;
  wire       [2:0]    resultStage_controlPipe_payload_twiceMode;
  wire                resultStage_controlPipe_payload_inpValidFlag;
  wire                resultStage_controlPipe_payload_oddValid;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rValid;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_frameStart;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_rowEnd;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_passMode;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_passValid;
  reg        [2:0]    diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_onceMode;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_onceValid;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_mainCompare;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_counterCompare;
  reg        [7:0]    diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_mainDiff;
  reg        [7:0]    diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_counterDiff;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_twiceCompValid;
  reg        [2:0]    diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_twiceMode;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_inpValidFlag;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_oddValid;
  wire                when_Stream_l368_31;
  wire                resultStage_pixelStream_valid;
  wire                resultStage_pixelStream_ready;
  reg        [7:0]    resultStage_pixelStream_payload;
  wire                when_SuperResolutionPart2_l451;
  wire                when_SuperResolutionPart2_l455;
  wire                when_SuperResolutionPart2_l459;
  wire                when_SuperResolutionPart2_l463;
  wire                when_SuperResolutionPart2_l474;
  wire                when_SuperResolutionPart2_l477;
  wire                when_SuperResolutionPart2_l482;
  wire                when_SuperResolutionPart2_l485;
  wire                when_SuperResolutionPart2_l491;
  wire                when_SuperResolutionPart2_l496;
  wire                resultStage_pixelStream_s2mPipe_valid;
  reg                 resultStage_pixelStream_s2mPipe_ready;
  wire       [7:0]    resultStage_pixelStream_s2mPipe_payload;
  reg                 resultStage_pixelStream_rValid;
  reg        [7:0]    resultStage_pixelStream_rData;
  wire                resultStage_resultStream_valid;
  wire                resultStage_resultStream_ready;
  wire       [7:0]    resultStage_resultStream_payload;
  reg                 resultStage_pixelStream_s2mPipe_rValid;
  reg        [7:0]    resultStage_pixelStream_s2mPipe_rData;
  wire                when_Stream_l368_32;
  wire                CICC1851_resultStage_mainOnePixelStream_ready;
  reg                 CICC1851_resultStage_mainOnePixelStream_ready_1;
  wire                CICC1851_resultStage_mainOnePixelStream_ready_2;
  wire                when_Stream_l438;
  reg                 resultsJoin_valid;
  wire                resultsJoin_ready;
  wire                pixelsStream_valid;
  wire                pixelsStream_ready;
  wire       [7:0]    pixelsStream_payload_pixel;
  wire                pixelsStream_payload_frameStart;
  wire                pixelsStream_payload_rowEnd;
  wire                pixelsStream_payload_inpValid;
  wire                pixelsStream_s2mPipe_valid;
  reg                 pixelsStream_s2mPipe_ready;
  wire       [7:0]    pixelsStream_s2mPipe_payload_pixel;
  wire                pixelsStream_s2mPipe_payload_frameStart;
  wire                pixelsStream_s2mPipe_payload_rowEnd;
  wire                pixelsStream_s2mPipe_payload_inpValid;
  reg                 pixelsStream_rValid;
  reg        [7:0]    pixelsStream_rData_pixel;
  reg                 pixelsStream_rData_frameStart;
  reg                 pixelsStream_rData_rowEnd;
  reg                 pixelsStream_rData_inpValid;
  wire                pixelsStream_s2mPipe_m2sPipe_valid;
  wire                pixelsStream_s2mPipe_m2sPipe_ready;
  wire       [7:0]    pixelsStream_s2mPipe_m2sPipe_payload_pixel;
  wire                pixelsStream_s2mPipe_m2sPipe_payload_frameStart;
  wire                pixelsStream_s2mPipe_m2sPipe_payload_rowEnd;
  wire                pixelsStream_s2mPipe_m2sPipe_payload_inpValid;
  reg                 pixelsStream_s2mPipe_rValid;
  reg        [7:0]    pixelsStream_s2mPipe_rData_pixel;
  reg                 pixelsStream_s2mPipe_rData_frameStart;
  reg                 pixelsStream_s2mPipe_rData_rowEnd;
  reg                 pixelsStream_s2mPipe_rData_inpValid;
  wire                when_Stream_l368_33;
  wire                controlStateMachine_wantExit;
  reg                 controlStateMachine_wantStart;
  wire                controlStateMachine_wantKill;
  wire                when_SuperResolutionPart2_l761;
  wire                controlStream_fire_4;
  wire                when_SuperResolutionPart2_l763;
  wire                controlStream_fire_5;
  wire                when_SuperResolutionPart2_l764;
  wire                controlStream_fire_6;
  wire                when_SuperResolutionPart2_l766;
  wire                controlStream_fire_7;
  wire                when_SuperResolutionPart2_l783;
  wire                when_SuperResolutionPart2_l785;
  wire                when_SuperResolutionPart2_l787;
  wire                when_SuperResolutionPart2_l789;
  wire                when_SuperResolutionPart2_l793;
  wire                when_SuperResolutionPart2_l796;
  wire                when_SuperResolutionPart2_l799;
  wire                when_SuperResolutionPart2_l802;
  reg        [2:0]    controlStateMachine_stateReg;
  reg        [2:0]    controlStateMachine_stateNext;
  wire                passPixels_fire_13;
  wire                passPixels_fire_14;
  wire                passPixels_fire_15;
  wire                passPixels_fire_16;
  wire                when_SuperResolutionPart2_l560;
  wire                controlStream_fire_8;
  wire                passPixels_fire_17;
  wire                when_SuperResolutionPart2_l573;
  wire                passPixels_fire_18;
  wire                when_SuperResolutionPart2_l578;
  wire                when_SuperResolutionPart2_l585;
  wire                when_SuperResolutionPart2_l588;
  wire                passPixels_fire_19;
  wire                when_SuperResolutionPart2_l590;
  wire                when_SuperResolutionPart2_l602;
  wire                when_SuperResolutionPart2_l603;
  wire                when_SuperResolutionPart2_l605;
  wire                when_SuperResolutionPart2_l606;
  wire                when_SuperResolutionPart2_l609;
  wire                controlStream_fire_9;
  wire                when_SuperResolutionPart2_l630;
  wire                controlStream_fire_10;
  wire                passPixels_fire_20;
  wire                when_SuperResolutionPart2_l642;
  wire                passPixels_fire_21;
  wire                when_SuperResolutionPart2_l647;
  wire                passPixels_fire_22;
  wire                when_SuperResolutionPart2_l653;
  wire                passPixels_fire_23;
  wire                when_SuperResolutionPart2_l662;
  wire                when_SuperResolutionPart2_l667;
  wire                when_SuperResolutionPart2_l668;
  wire                controlStream_fire_11;
  `ifndef SYNTHESIS
  reg [39:0] controlStateMachine_stateReg_string;
  reg [39:0] controlStateMachine_stateNext_string;
  `endif

  reg [7:0] lineBufferOne [0:1919];
  reg [7:0] lineBufferTwo [0:1919];
  reg [7:0] lineBufferOdd [0:1919];

  assign CICC1851_bufferRowCount_valueNext_1 = bufferRowCount_willIncrement;
  assign CICC1851_bufferRowCount_valueNext = {10'd0, CICC1851_bufferRowCount_valueNext_1};
  assign CICC1851_bufferWAddr_valueNext_1 = bufferWAddr_willIncrement;
  assign CICC1851_bufferWAddr_valueNext = {10'd0, CICC1851_bufferWAddr_valueNext_1};
  assign CICC1851_outPixelAddr_valueNext_1 = outPixelAddr_willIncrement;
  assign CICC1851_outPixelAddr_valueNext = {11'd0, CICC1851_outPixelAddr_valueNext_1};
  assign CICC1851_outRowCount_valueNext_1 = outRowCount_willIncrement;
  assign CICC1851_outRowCount_valueNext = {11'd0, CICC1851_outRowCount_valueNext_1};
  assign CICC1851_alreadySendRow_valueNext_1 = alreadySendRow_willIncrement;
  assign CICC1851_alreadySendRow_valueNext = {11'd0, CICC1851_alreadySendRow_valueNext_1};
  assign CICC1851_alreadySendCountInRow_valueNext_1 = alreadySendCountInRow_willIncrement;
  assign CICC1851_alreadySendCountInRow_valueNext = {11'd0, CICC1851_alreadySendCountInRow_valueNext_1};
  assign CICC1851_mainAddrOne = (outPixelAddr_value / 2'b10);
  assign CICC1851_counterAddrOne = (outPixelAddr_value / 2'b10);
  assign CICC1851_mainAddrTwo = (outPixelAddr_value / 2'b10);
  assign CICC1851_counterAddrTwo = (outPixelAddr_value / 2'b10);
  assign CICC1851_oddAddr = (outPixelAddr_value / 2'b10);
  assign CICC1851_when_SuperResolutionPart2_l181 = {1'd0, bufferWAddr_value};
  assign CICC1851_when_SuperResolutionPart2_l181_1 = (CICC1851_when_SuperResolutionPart2_l181_2 - 12'h002);
  assign CICC1851_when_SuperResolutionPart2_l181_2 = (2'b10 * bmpWidth);
  assign CICC1851_when_SuperResolutionPart2_l182 = {1'd0, bufferRowCount_value};
  assign CICC1851_when_SuperResolutionPart2_l182_1 = (CICC1851_when_SuperResolutionPart2_l182_2 - 12'h002);
  assign CICC1851_when_SuperResolutionPart2_l182_2 = (2'b10 * bmpHeight);
  assign CICC1851_when_SuperResolutionPart2_l195 = (bufferRowCount_value % 2'b10);
  assign CICC1851_when_SuperResolutionPart2_l218 = (outRowCount_value % 3'b100);
  assign CICC1851_when_SuperResolutionPart2_l234 = {1'd0, alreadySendCountInRow_value};
  assign CICC1851_when_SuperResolutionPart2_l234_1 = (CICC1851_when_SuperResolutionPart2_l234_2 - 13'h0002);
  assign CICC1851_when_SuperResolutionPart2_l234_2 = (3'b100 * bmpWidth);
  assign CICC1851_when_SuperResolutionPart2_l235 = {1'd0, alreadySendRow_value};
  assign CICC1851_when_SuperResolutionPart2_l235_1 = (CICC1851_when_SuperResolutionPart2_l235_2 - 13'h0002);
  assign CICC1851_when_SuperResolutionPart2_l235_2 = (3'b100 * bmpHeight);
  assign CICC1851_resultStage_pixelStream_payload = (CICC1851_resultStage_pixelStream_payload_1 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_1 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_2 = (CICC1851_resultStage_pixelStream_payload_3 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_3 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_4 = (CICC1851_resultStage_pixelStream_payload_5 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_5 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_mainTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_6 = (CICC1851_resultStage_pixelStream_payload_7 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_7 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_mainOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_8 = (CICC1851_resultStage_pixelStream_payload_9 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_9 = ({1'b0,diffStage_counterOnePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_10 = (CICC1851_resultStage_pixelStream_payload_11 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_11 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_mainTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_12 = (CICC1851_resultStage_pixelStream_payload_13 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_13 = ({1'b0,diffStage_counterOnePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_14 = (CICC1851_resultStage_pixelStream_payload_15 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_15 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_mainTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_16 = (CICC1851_resultStage_pixelStream_payload_17 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_17 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_18 = (CICC1851_resultStage_pixelStream_payload_19 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_19 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_when_SuperResolutionPart2_l763 = {1'd0, outPixelAddr_value};
  assign CICC1851_when_SuperResolutionPart2_l763_1 = (CICC1851_when_SuperResolutionPart2_l763_2 - 13'h0002);
  assign CICC1851_when_SuperResolutionPart2_l763_2 = (3'b100 * bmpWidth);
  assign CICC1851_when_SuperResolutionPart2_l764 = {1'd0, outRowCount_value};
  assign CICC1851_when_SuperResolutionPart2_l764_1 = (CICC1851_when_SuperResolutionPart2_l764_2 - 13'h0002);
  assign CICC1851_when_SuperResolutionPart2_l764_2 = (3'b100 * bmpHeight);
  assign CICC1851_when_SuperResolutionPart2_l783 = (outRowCount_value % 3'b100);
  assign CICC1851_when_SuperResolutionPart2_l785 = (outRowCount_value % 3'b100);
  assign CICC1851_when_SuperResolutionPart2_l787 = (outRowCount_value % 3'b100);
  assign CICC1851_when_SuperResolutionPart2_l789 = (outRowCount_value % 3'b100);
  assign CICC1851_when_SuperResolutionPart2_l793 = (outPixelAddr_value % 3'b100);
  assign CICC1851_when_SuperResolutionPart2_l796 = (outPixelAddr_value % 3'b100);
  assign CICC1851_when_SuperResolutionPart2_l799 = (outPixelAddr_value % 3'b100);
  assign CICC1851_when_SuperResolutionPart2_l802 = (outPixelAddr_value % 3'b100);
  assign CICC1851_when_SuperResolutionPart2_l560 = (2'b10 * bufferWAddr_value);
  assign CICC1851_when_SuperResolutionPart2_l560_1 = {1'd0, outPixelAddr_value};
  assign CICC1851_when_SuperResolutionPart2_l602 = (2'b10 * bufferWAddr_value);
  assign CICC1851_when_SuperResolutionPart2_l602_1 = (CICC1851_when_SuperResolutionPart2_l602_2 + {1'b0,outPixelAddr_value});
  assign CICC1851_when_SuperResolutionPart2_l602_3 = {1'b0,2'b10};
  assign CICC1851_when_SuperResolutionPart2_l602_2 = {10'd0, CICC1851_when_SuperResolutionPart2_l602_3};
  assign CICC1851_when_SuperResolutionPart2_l603 = (2'b10 * bufferWAddr_value);
  assign CICC1851_when_SuperResolutionPart2_l603_1 = {1'd0, outPixelAddr_value};
  assign CICC1851_when_SuperResolutionPart2_l605 = (2'b10 * bufferWAddr_value);
  assign CICC1851_when_SuperResolutionPart2_l605_1 = (CICC1851_when_SuperResolutionPart2_l605_2 + {1'b0,outPixelAddr_value});
  assign CICC1851_when_SuperResolutionPart2_l605_3 = {1'b0,2'b11};
  assign CICC1851_when_SuperResolutionPart2_l605_2 = {10'd0, CICC1851_when_SuperResolutionPart2_l605_3};
  assign CICC1851_when_SuperResolutionPart2_l606 = (2'b10 * bufferWAddr_value);
  assign CICC1851_when_SuperResolutionPart2_l606_1 = (CICC1851_when_SuperResolutionPart2_l606_2 + {1'b0,outPixelAddr_value});
  assign CICC1851_when_SuperResolutionPart2_l606_3 = {1'b0,1'b1};
  assign CICC1851_when_SuperResolutionPart2_l606_2 = {11'd0, CICC1851_when_SuperResolutionPart2_l606_3};
  assign CICC1851_when_SuperResolutionPart2_l609 = (outPixelAddr_value % 2'b10);
  assign CICC1851_mainAddrOne_1 = (CICC1851_mainAddrOne_2 / 2'b10);
  assign CICC1851_mainAddrOne_2 = (outPixelAddr_value - 12'h002);
  assign CICC1851_mainAddrTwo_1 = (CICC1851_mainAddrTwo_2 / 2'b10);
  assign CICC1851_mainAddrTwo_2 = (outPixelAddr_value - 12'h002);
  assign CICC1851_when_SuperResolutionPart2_l667 = (CICC1851_when_SuperResolutionPart2_l667_1 - 13'h0002);
  assign CICC1851_when_SuperResolutionPart2_l667_1 = (2'b10 * bufferWAddr_value);
  assign CICC1851_when_SuperResolutionPart2_l667_2 = (CICC1851_when_SuperResolutionPart2_l667_3 + {1'b0,outPixelAddr_value});
  assign CICC1851_when_SuperResolutionPart2_l667_4 = {1'b0,1'b1};
  assign CICC1851_when_SuperResolutionPart2_l667_3 = {11'd0, CICC1851_when_SuperResolutionPart2_l667_4};
  assign CICC1851_when_SuperResolutionPart2_l668 = (2'b10 * bufferWAddr_value);
  assign CICC1851_when_SuperResolutionPart2_l668_1 = (CICC1851_when_SuperResolutionPart2_l668_2 + {1'b0,outPixelAddr_value});
  assign CICC1851_when_SuperResolutionPart2_l668_3 = {1'b0,1'b1};
  assign CICC1851_when_SuperResolutionPart2_l668_2 = {11'd0, CICC1851_when_SuperResolutionPart2_l668_3};
  assign CICC1851_mainAddrOne_3 = (CICC1851_mainAddrOne_4 / 2'b10);
  assign CICC1851_mainAddrOne_4 = (outPixelAddr_value - 12'h002);
  assign CICC1851_mainAddrTwo_3 = (CICC1851_mainAddrTwo_4 / 2'b10);
  assign CICC1851_mainAddrTwo_4 = (outPixelAddr_value - 12'h002);
  assign CICC1851_controls_onceMode = 2'b10;
  assign CICC1851_controls_onceMode_1 = 2'b11;
  assign CICC1851_mainAddrOne_5 = (CICC1851_mainAddrOne_6 / 2'b10);
  assign CICC1851_mainAddrOne_6 = (outPixelAddr_value - 12'h003);
  assign CICC1851_counterAddrOne_1 = (CICC1851_counterAddrOne_2 / 2'b10);
  assign CICC1851_counterAddrOne_2 = (outPixelAddr_value - 12'h003);
  assign CICC1851_counterAddrOne_3 = (CICC1851_counterAddrOne_4 / 2'b10);
  assign CICC1851_counterAddrOne_4 = (12'h001 + outPixelAddr_value);
  assign CICC1851_controls_onceMode_2 = 1'b1;
  assign CICC1851_mainAddrTwo_5 = (CICC1851_mainAddrTwo_6 / 2'b10);
  assign CICC1851_mainAddrTwo_6 = (outPixelAddr_value - 12'h003);
  assign CICC1851_counterAddrTwo_1 = (CICC1851_counterAddrTwo_2 / 2'b10);
  assign CICC1851_counterAddrTwo_2 = (outPixelAddr_value - 12'h003);
  assign CICC1851_counterAddrTwo_3 = (CICC1851_counterAddrTwo_4 / 2'b10);
  assign CICC1851_counterAddrTwo_4 = (12'h001 + outPixelAddr_value);
  assign CICC1851_mainAddrOne_7 = (CICC1851_mainAddrOne_8 / 2'b10);
  assign CICC1851_mainAddrOne_8 = (outPixelAddr_value - 12'h003);
  assign CICC1851_mainAddrOne_9 = (CICC1851_mainAddrOne_10 / 2'b10);
  assign CICC1851_mainAddrOne_10 = (outPixelAddr_value - 12'h003);
  assign CICC1851_counterAddrOne_5 = (CICC1851_counterAddrOne_6 / 2'b10);
  assign CICC1851_counterAddrOne_6 = (CICC1851_counterAddrOne_7 + {1'b0,outPixelAddr_value});
  assign CICC1851_counterAddrOne_8 = {1'b0,1'b1};
  assign CICC1851_counterAddrOne_7 = {11'd0, CICC1851_counterAddrOne_8};
  assign CICC1851_controls_twiceMode = 2'b10;
  assign CICC1851_mainAddrTwo_7 = (CICC1851_mainAddrTwo_8 / 2'b10);
  assign CICC1851_mainAddrTwo_8 = (outPixelAddr_value - 12'h003);
  assign CICC1851_controls_twiceMode_1 = 2'b11;
  assign CICC1851_mainAddrTwo_9 = (CICC1851_mainAddrTwo_10 / 2'b10);
  assign CICC1851_mainAddrTwo_10 = (outPixelAddr_value - 12'h003);
  assign CICC1851_counterAddrTwo_5 = (CICC1851_counterAddrTwo_6 / 2'b10);
  assign CICC1851_counterAddrTwo_6 = (CICC1851_counterAddrTwo_7 + {1'b0,outPixelAddr_value});
  assign CICC1851_counterAddrTwo_8 = {1'b0,1'b1};
  assign CICC1851_counterAddrTwo_7 = {11'd0, CICC1851_counterAddrTwo_8};
  assign CICC1851_mainAddrOne_11 = (CICC1851_mainAddrOne_12 / 2'b10);
  assign CICC1851_mainAddrOne_12 = (outPixelAddr_value - 12'h003);
  assign CICC1851_counterAddrTwo_9 = (CICC1851_counterAddrTwo_10 / 2'b10);
  assign CICC1851_counterAddrTwo_10 = (outPixelAddr_value - 12'h003);
  assign CICC1851_mainAddrTwo_11 = (CICC1851_mainAddrTwo_12 / 2'b10);
  assign CICC1851_mainAddrTwo_12 = (outPixelAddr_value - 12'h003);
  assign CICC1851_counterAddrOne_9 = (CICC1851_counterAddrOne_10 / 2'b10);
  assign CICC1851_counterAddrOne_10 = (outPixelAddr_value - 12'h003);
  assign CICC1851_mainAddrTwo_13 = (CICC1851_mainAddrTwo_14 / 2'b10);
  assign CICC1851_mainAddrTwo_14 = ({1'b0,outPixelAddr_value} + CICC1851_mainAddrTwo_15);
  assign CICC1851_mainAddrTwo_16 = {1'b0,1'b1};
  assign CICC1851_mainAddrTwo_15 = {11'd0, CICC1851_mainAddrTwo_16};
  assign CICC1851_counterAddrOne_11 = (CICC1851_counterAddrOne_12 / 2'b10);
  assign CICC1851_counterAddrOne_12 = ({1'b0,outPixelAddr_value} + CICC1851_counterAddrOne_13);
  assign CICC1851_counterAddrOne_14 = {1'b0,1'b1};
  assign CICC1851_counterAddrOne_13 = {11'd0, CICC1851_counterAddrOne_14};
  assign CICC1851_controls_twiceMode_2 = 1'b1;
  assign CICC1851_mainAddrTwo_17 = (CICC1851_mainAddrTwo_18 / 2'b10);
  assign CICC1851_mainAddrTwo_18 = (outPixelAddr_value - 12'h003);
  assign CICC1851_counterAddrOne_15 = (CICC1851_counterAddrOne_16 / 2'b10);
  assign CICC1851_counterAddrOne_16 = (outPixelAddr_value - 12'h003);
  assign CICC1851_mainAddrOne_13 = (CICC1851_mainAddrOne_14 / 2'b10);
  assign CICC1851_mainAddrOne_14 = (outPixelAddr_value - 12'h003);
  assign CICC1851_counterAddrTwo_11 = (CICC1851_counterAddrTwo_12 / 2'b10);
  assign CICC1851_counterAddrTwo_12 = (outPixelAddr_value - 12'h003);
  assign CICC1851_mainAddrOne_15 = (CICC1851_mainAddrOne_16 / 2'b10);
  assign CICC1851_mainAddrOne_16 = ({1'b0,outPixelAddr_value} + CICC1851_mainAddrOne_17);
  assign CICC1851_mainAddrOne_18 = {1'b0,1'b1};
  assign CICC1851_mainAddrOne_17 = {11'd0, CICC1851_mainAddrOne_18};
  assign CICC1851_counterAddrTwo_13 = (CICC1851_counterAddrTwo_14 / 2'b10);
  assign CICC1851_counterAddrTwo_14 = ({1'b0,outPixelAddr_value} + CICC1851_counterAddrTwo_15);
  assign CICC1851_counterAddrTwo_16 = {1'b0,1'b1};
  assign CICC1851_counterAddrTwo_15 = {11'd0, CICC1851_counterAddrTwo_16};
  assign CICC1851_lineBufferOne_port = passPixels_payload_pixel;
  assign CICC1851_lineBufferOne_port_1 = (passPixels_fire_6 && (bufferSwitch == 2'b00));
  assign CICC1851_lineBufferTwo_port = passPixels_payload_pixel;
  assign CICC1851_lineBufferTwo_port_1 = (passPixels_fire_8 && (bufferSwitch == 2'b10));
  assign CICC1851_lineBufferOdd_port = passPixels_payload_pixel;
  assign CICC1851_lineBufferOdd_port_1 = (passPixels_fire_7 && (bufferSwitch == 2'b01));
  always @(posedge clk) begin
    if(CICC1851_lineBufferOne_port_1) begin
      lineBufferOne[bufferWAddr_value] <= CICC1851_lineBufferOne_port;
    end
  end

  always @(posedge clk) begin
    if(mainAddrOneStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferOne_port1 <= lineBufferOne[mainAddrOneStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(counterAddrOneStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferOne_port2 <= lineBufferOne[counterAddrOneStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(CICC1851_lineBufferTwo_port_1) begin
      lineBufferTwo[bufferWAddr_value] <= CICC1851_lineBufferTwo_port;
    end
  end

  always @(posedge clk) begin
    if(mainAddrTwoStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferTwo_port1 <= lineBufferTwo[mainAddrTwoStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(counterAddrTwoStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferTwo_port2 <= lineBufferTwo[counterAddrTwoStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(CICC1851_lineBufferOdd_port_1) begin
      lineBufferOdd[bufferWAddr_value] <= CICC1851_lineBufferOdd_port;
    end
  end

  always @(posedge clk) begin
    if(oddAddrStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferOdd_port1 <= lineBufferOdd[oddAddrStream_s2mPipe_m2sPipe_payload];
    end
  end

  StreamFork_2 diffStage_controlPipe_fork (
    .io_input_valid                      (diffStage_controlPipe_valid                                     ), //i
    .io_input_ready                      (diffStage_controlPipe_fork_io_input_ready                       ), //o
    .io_input_payload_frameStart         (diffStage_controlPipe_payload_frameStart                        ), //i
    .io_input_payload_rowEnd             (diffStage_controlPipe_payload_rowEnd                            ), //i
    .io_input_payload_passMode           (diffStage_controlPipe_payload_passMode                          ), //i
    .io_input_payload_passValid          (diffStage_controlPipe_payload_passValid                         ), //i
    .io_input_payload_onceMode           (diffStage_controlPipe_payload_onceMode[2:0]                     ), //i
    .io_input_payload_onceValid          (diffStage_controlPipe_payload_onceValid                         ), //i
    .io_input_payload_mainCompare        (diffStage_controlPipe_payload_mainCompare                       ), //i
    .io_input_payload_counterCompare     (diffStage_controlPipe_payload_counterCompare                    ), //i
    .io_input_payload_mainDiff           (diffStage_controlPipe_payload_mainDiff[7:0]                     ), //i
    .io_input_payload_counterDiff        (diffStage_controlPipe_payload_counterDiff[7:0]                  ), //i
    .io_input_payload_twiceCompValid     (diffStage_controlPipe_payload_twiceCompValid                    ), //i
    .io_input_payload_twiceMode          (diffStage_controlPipe_payload_twiceMode[2:0]                    ), //i
    .io_input_payload_inpValidFlag       (diffStage_controlPipe_payload_inpValidFlag                      ), //i
    .io_input_payload_oddValid           (diffStage_controlPipe_payload_oddValid                          ), //i
    .io_outputs_0_valid                  (diffStage_controlPipe_fork_io_outputs_0_valid                   ), //o
    .io_outputs_0_ready                  (diffStage_controlPipe_fork_io_outputs_0_translated_ready        ), //i
    .io_outputs_0_payload_frameStart     (diffStage_controlPipe_fork_io_outputs_0_payload_frameStart      ), //o
    .io_outputs_0_payload_rowEnd         (diffStage_controlPipe_fork_io_outputs_0_payload_rowEnd          ), //o
    .io_outputs_0_payload_passMode       (diffStage_controlPipe_fork_io_outputs_0_payload_passMode        ), //o
    .io_outputs_0_payload_passValid      (diffStage_controlPipe_fork_io_outputs_0_payload_passValid       ), //o
    .io_outputs_0_payload_onceMode       (diffStage_controlPipe_fork_io_outputs_0_payload_onceMode[2:0]   ), //o
    .io_outputs_0_payload_onceValid      (diffStage_controlPipe_fork_io_outputs_0_payload_onceValid       ), //o
    .io_outputs_0_payload_mainCompare    (diffStage_controlPipe_fork_io_outputs_0_payload_mainCompare     ), //o
    .io_outputs_0_payload_counterCompare (diffStage_controlPipe_fork_io_outputs_0_payload_counterCompare  ), //o
    .io_outputs_0_payload_mainDiff       (diffStage_controlPipe_fork_io_outputs_0_payload_mainDiff[7:0]   ), //o
    .io_outputs_0_payload_counterDiff    (diffStage_controlPipe_fork_io_outputs_0_payload_counterDiff[7:0]), //o
    .io_outputs_0_payload_twiceCompValid (diffStage_controlPipe_fork_io_outputs_0_payload_twiceCompValid  ), //o
    .io_outputs_0_payload_twiceMode      (diffStage_controlPipe_fork_io_outputs_0_payload_twiceMode[2:0]  ), //o
    .io_outputs_0_payload_inpValidFlag   (diffStage_controlPipe_fork_io_outputs_0_payload_inpValidFlag    ), //o
    .io_outputs_0_payload_oddValid       (diffStage_controlPipe_fork_io_outputs_0_payload_oddValid        ), //o
    .io_outputs_1_valid                  (diffStage_controlPipe_fork_io_outputs_1_valid                   ), //o
    .io_outputs_1_ready                  (resultStage_pixelStream_ready                                   ), //i
    .io_outputs_1_payload_frameStart     (diffStage_controlPipe_fork_io_outputs_1_payload_frameStart      ), //o
    .io_outputs_1_payload_rowEnd         (diffStage_controlPipe_fork_io_outputs_1_payload_rowEnd          ), //o
    .io_outputs_1_payload_passMode       (diffStage_controlPipe_fork_io_outputs_1_payload_passMode        ), //o
    .io_outputs_1_payload_passValid      (diffStage_controlPipe_fork_io_outputs_1_payload_passValid       ), //o
    .io_outputs_1_payload_onceMode       (diffStage_controlPipe_fork_io_outputs_1_payload_onceMode[2:0]   ), //o
    .io_outputs_1_payload_onceValid      (diffStage_controlPipe_fork_io_outputs_1_payload_onceValid       ), //o
    .io_outputs_1_payload_mainCompare    (diffStage_controlPipe_fork_io_outputs_1_payload_mainCompare     ), //o
    .io_outputs_1_payload_counterCompare (diffStage_controlPipe_fork_io_outputs_1_payload_counterCompare  ), //o
    .io_outputs_1_payload_mainDiff       (diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff[7:0]   ), //o
    .io_outputs_1_payload_counterDiff    (diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff[7:0]), //o
    .io_outputs_1_payload_twiceCompValid (diffStage_controlPipe_fork_io_outputs_1_payload_twiceCompValid  ), //o
    .io_outputs_1_payload_twiceMode      (diffStage_controlPipe_fork_io_outputs_1_payload_twiceMode[2:0]  ), //o
    .io_outputs_1_payload_inpValidFlag   (diffStage_controlPipe_fork_io_outputs_1_payload_inpValidFlag    ), //o
    .io_outputs_1_payload_oddValid       (diffStage_controlPipe_fork_io_outputs_1_payload_oddValid        )  //o
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_4_BOOT : controlStateMachine_stateReg_string = "BOOT ";
      controlStateMachine_enumDef_4_HOLD : controlStateMachine_stateReg_string = "HOLD ";
      controlStateMachine_enumDef_4_PASS : controlStateMachine_stateReg_string = "PASS ";
      controlStateMachine_enumDef_4_ONCE : controlStateMachine_stateReg_string = "ONCE ";
      controlStateMachine_enumDef_4_TWICE : controlStateMachine_stateReg_string = "TWICE";
      default : controlStateMachine_stateReg_string = "?????";
    endcase
  end
  always @(*) begin
    case(controlStateMachine_stateNext)
      controlStateMachine_enumDef_4_BOOT : controlStateMachine_stateNext_string = "BOOT ";
      controlStateMachine_enumDef_4_HOLD : controlStateMachine_stateNext_string = "HOLD ";
      controlStateMachine_enumDef_4_PASS : controlStateMachine_stateNext_string = "PASS ";
      controlStateMachine_enumDef_4_ONCE : controlStateMachine_stateNext_string = "ONCE ";
      controlStateMachine_enumDef_4_TWICE : controlStateMachine_stateNext_string = "TWICE";
      default : controlStateMachine_stateNext_string = "?????";
    endcase
  end
  `endif

  always @(*) begin
    pixelsIn_ready = 1'b0;
    pixelsIn_ready = (! pixelsIn_rValid);
  end

  always @(*) begin
    pixelsOut_valid = 1'b0;
    pixelsOut_valid = pixelsStream_s2mPipe_m2sPipe_valid;
  end

  always @(*) begin
    pixelsOut_payload_pixel = 8'h0;
    pixelsOut_payload_pixel = pixelsStream_s2mPipe_m2sPipe_payload_pixel;
  end

  always @(*) begin
    pixelsOut_payload_frameStart = 1'b0;
    pixelsOut_payload_frameStart = pixelsStream_s2mPipe_m2sPipe_payload_frameStart;
  end

  always @(*) begin
    pixelsOut_payload_rowEnd = 1'b0;
    pixelsOut_payload_rowEnd = pixelsStream_s2mPipe_m2sPipe_payload_rowEnd;
  end

  always @(*) begin
    pixelsOut_payload_inpValid = 1'b0;
    pixelsOut_payload_inpValid = pixelsStream_s2mPipe_m2sPipe_payload_inpValid;
  end

  always @(*) begin
    startOut = 1'b0;
    startOut = slaveStart;
  end

  always @(*) begin
    inpTwoDoneOut = 1'b0;
    inpTwoDoneOut = inpTwoDone;
  end

  assign when_SuperResolutionPart2_l40 = (inpThreeDoneIn || (startIn && (! startIn_regNext)));
  assign when_SuperResolutionPart2_l43 = (! startIn);
  assign when_SuperResolutionPart2_l46 = (startIn && (! readDone));
  assign when_SuperResolutionPart2_l46_1 = (! startIn);
  assign pixelsIn_fire = (pixelsIn_valid && pixelsIn_ready);
  assign when_SuperResolutionPart2_l49 = ((! inpThreeDoneIn) && pixelsIn_fire);
  assign when_SuperResolutionPart2_l49_1 = (inpThreeDoneIn || (! startIn));
  assign when_SuperResolutionPart2_l64 = (! startIn);
  assign when_SuperResolutionPart2_l67 = (! startIn);
  always @(*) begin
    bufferRowCount_willIncrement = 1'b0;
    if(when_SuperResolutionPart2_l185) begin
      if(!bufferReachFinalRow) begin
        bufferRowCount_willIncrement = 1'b1;
      end
    end
  end

  always @(*) begin
    bufferRowCount_willClear = 1'b0;
    if(when_SuperResolutionPart2_l185) begin
      if(bufferReachFinalRow) begin
        bufferRowCount_willClear = 1'b1;
      end
    end
  end

  assign bufferRowCount_willOverflowIfInc = (bufferRowCount_value == 11'h438);
  assign bufferRowCount_willOverflow = (bufferRowCount_willOverflowIfInc && bufferRowCount_willIncrement);
  always @(*) begin
    if(bufferRowCount_willOverflow) begin
      bufferRowCount_valueNext = 11'h0;
    end else begin
      bufferRowCount_valueNext = (bufferRowCount_value + CICC1851_bufferRowCount_valueNext);
    end
    if(bufferRowCount_willClear) begin
      bufferRowCount_valueNext = 11'h0;
    end
  end

  assign when_SuperResolutionPart2_l76 = ((startIn && (! holdBuffer)) && (! writeDone));
  assign when_SuperResolutionPart2_l76_1 = (((! startIn) || holdBuffer) || writeDone);
  assign when_SuperResolutionPart2_l82 = (! startRead);
  always @(*) begin
    bufferWAddr_willIncrement = 1'b0;
    if(passPixels_fire_9) begin
      if(!passPixels_payload_rowEnd) begin
        bufferWAddr_willIncrement = 1'b1;
      end
    end
  end

  always @(*) begin
    bufferWAddr_willClear = 1'b0;
    if(passPixels_fire_9) begin
      if(passPixels_payload_rowEnd) begin
        bufferWAddr_willClear = 1'b1;
      end
    end
  end

  assign bufferWAddr_willOverflowIfInc = (bufferWAddr_value == 11'h77f);
  assign bufferWAddr_willOverflow = (bufferWAddr_willOverflowIfInc && bufferWAddr_willIncrement);
  always @(*) begin
    if(bufferWAddr_willOverflow) begin
      bufferWAddr_valueNext = 11'h0;
    end else begin
      bufferWAddr_valueNext = (bufferWAddr_value + CICC1851_bufferWAddr_valueNext);
    end
    if(bufferWAddr_willClear) begin
      bufferWAddr_valueNext = 11'h0;
    end
  end

  always @(*) begin
    outPixelAddr_willIncrement = 1'b0;
    if(when_SuperResolutionPart2_l761) begin
      if(controlStream_fire_7) begin
        if(!outReachRowEnd) begin
          outPixelAddr_willIncrement = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    outPixelAddr_willClear = 1'b0;
    if(when_SuperResolutionPart2_l761) begin
      if(controlStream_fire_7) begin
        if(outReachRowEnd) begin
          outPixelAddr_willClear = 1'b1;
        end
      end
    end
  end

  assign outPixelAddr_willOverflowIfInc = (outPixelAddr_value == 12'heff);
  assign outPixelAddr_willOverflow = (outPixelAddr_willOverflowIfInc && outPixelAddr_willIncrement);
  always @(*) begin
    if(outPixelAddr_willOverflow) begin
      outPixelAddr_valueNext = 12'h0;
    end else begin
      outPixelAddr_valueNext = (outPixelAddr_value + CICC1851_outPixelAddr_valueNext);
    end
    if(outPixelAddr_willClear) begin
      outPixelAddr_valueNext = 12'h0;
    end
  end

  always @(*) begin
    outRowCount_willIncrement = 1'b0;
    if(when_SuperResolutionPart2_l761) begin
      if(when_SuperResolutionPart2_l766) begin
        if(!outReachFinalRow) begin
          outRowCount_willIncrement = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    outRowCount_willClear = 1'b0;
    if(when_SuperResolutionPart2_l761) begin
      if(when_SuperResolutionPart2_l766) begin
        if(outReachFinalRow) begin
          outRowCount_willClear = 1'b1;
        end
      end
    end
  end

  assign outRowCount_willOverflowIfInc = (outRowCount_value == 12'h870);
  assign outRowCount_willOverflow = (outRowCount_willOverflowIfInc && outRowCount_willIncrement);
  always @(*) begin
    if(outRowCount_willOverflow) begin
      outRowCount_valueNext = 12'h0;
    end else begin
      outRowCount_valueNext = (outRowCount_value + CICC1851_outRowCount_valueNext);
    end
    if(outRowCount_willClear) begin
      outRowCount_valueNext = 12'h0;
    end
  end

  always @(*) begin
    alreadySendRow_willIncrement = 1'b0;
    if(pixelsOut_fire_2) begin
      if(alreadyReachRowEnd) begin
        if(!alreadyReachFinalRow) begin
          alreadySendRow_willIncrement = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    alreadySendRow_willClear = 1'b0;
    if(pixelsOut_fire_2) begin
      if(alreadyReachRowEnd) begin
        if(alreadyReachFinalRow) begin
          alreadySendRow_willClear = 1'b1;
        end
      end
    end
  end

  assign alreadySendRow_willOverflowIfInc = (alreadySendRow_value == 12'h870);
  assign alreadySendRow_willOverflow = (alreadySendRow_willOverflowIfInc && alreadySendRow_willIncrement);
  always @(*) begin
    if(alreadySendRow_willOverflow) begin
      alreadySendRow_valueNext = 12'h0;
    end else begin
      alreadySendRow_valueNext = (alreadySendRow_value + CICC1851_alreadySendRow_valueNext);
    end
    if(alreadySendRow_willClear) begin
      alreadySendRow_valueNext = 12'h0;
    end
  end

  always @(*) begin
    alreadySendCountInRow_willIncrement = 1'b0;
    if(pixelsOut_fire_2) begin
      if(!alreadyReachRowEnd) begin
        alreadySendCountInRow_willIncrement = 1'b1;
      end
    end
  end

  always @(*) begin
    alreadySendCountInRow_willClear = 1'b0;
    if(pixelsOut_fire_2) begin
      if(alreadyReachRowEnd) begin
        alreadySendCountInRow_willClear = 1'b1;
      end
    end
  end

  assign alreadySendCountInRow_willOverflowIfInc = (alreadySendCountInRow_value == 12'heff);
  assign alreadySendCountInRow_willOverflow = (alreadySendCountInRow_willOverflowIfInc && alreadySendCountInRow_willIncrement);
  always @(*) begin
    if(alreadySendCountInRow_willOverflow) begin
      alreadySendCountInRow_valueNext = 12'h0;
    end else begin
      alreadySendCountInRow_valueNext = (alreadySendCountInRow_value + CICC1851_alreadySendCountInRow_valueNext);
    end
    if(alreadySendCountInRow_willClear) begin
      alreadySendCountInRow_valueNext = 12'h0;
    end
  end

  assign when_SuperResolutionPart2_l106 = (((! startIn) && startIn_regNext_1) || inpTwoDone);
  assign when_SuperResolutionPart2_l108 = (((! startIn) && startIn_regNext_2) || inpTwoDone);
  assign when_SuperResolutionPart2_l109 = (((! startIn) && startIn_regNext_3) || inpTwoDone);
  assign when_SuperResolutionPart2_l110 = (((! startIn) && startIn_regNext_4) || inpTwoDone);
  assign when_SuperResolutionPart2_l111 = (((! startIn) && startIn_regNext_5) || inpTwoDone);
  assign when_SuperResolutionPart2_l113 = (((! startIn) && startIn_regNext_6) || inpTwoDone);
  assign when_SuperResolutionPart2_l114 = (((! startIn) && startIn_regNext_7) || inpTwoDone);
  assign when_SuperResolutionPart2_l115 = (((! startIn) && startIn_regNext_8) || inpTwoDone);
  assign when_SuperResolutionPart2_l116 = (((! startIn) && startIn_regNext_9) || inpTwoDone);
  assign when_SuperResolutionPart2_l120 = (((! startIn) && startIn_regNext_10) || inpTwoDone);
  assign when_SuperResolutionPart2_l121 = (((! startIn) && startIn_regNext_11) || inpTwoDone);
  assign when_SuperResolutionPart2_l122 = (((! startIn) && startIn_regNext_12) || inpTwoDone);
  assign when_SuperResolutionPart2_l123 = (((! startIn) && startIn_regNext_13) || inpTwoDone);
  assign when_SuperResolutionPart2_l124 = (((! startIn) && startIn_regNext_14) || inpTwoDone);
  assign when_SuperResolutionPart2_l125 = (((! startIn) && startIn_regNext_15) || inpTwoDone);
  assign when_SuperResolutionPart2_l126 = (((! startIn) && startIn_regNext_16) || inpTwoDone);
  assign when_SuperResolutionPart2_l134 = (! startRead);
  always @(*) begin
    mainAddrOne = CICC1851_mainAddrOne[10:0];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_4_HOLD : begin
      end
      controlStateMachine_enumDef_4_PASS : begin
        if(!twoInFourOutRow) begin
          if(oneInFourOutRow) begin
            if(nextRowBuffer) begin
              if(twoInFourOutPixelAddr) begin
                mainAddrOne = CICC1851_mainAddrOne_1[10:0];
              end
            end
          end
        end
      end
      controlStateMachine_enumDef_4_ONCE : begin
        if(threeInFourOutRow) begin
          if(twoInFourOutPixelAddr) begin
            mainAddrOne = CICC1851_mainAddrOne_3[10:0];
          end
        end else begin
          if(nextRowBuffer) begin
            mainAddrOne = CICC1851_mainAddrOne_5[10:0];
          end
        end
      end
      controlStateMachine_enumDef_4_TWICE : begin
        if(outReachFinalRow) begin
          if(nextRowBuffer) begin
            if(outReachRowEnd) begin
              mainAddrOne = CICC1851_mainAddrOne_7[10:0];
            end else begin
              mainAddrOne = CICC1851_mainAddrOne_9[10:0];
            end
          end
        end else begin
          if(nextRowBuffer) begin
            mainAddrOne = CICC1851_mainAddrOne_11[10:0];
          end else begin
            if(outReachRowEnd) begin
              mainAddrOne = CICC1851_mainAddrOne_13[10:0];
            end else begin
              mainAddrOne = CICC1851_mainAddrOne_15[10:0];
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    counterAddrOne = CICC1851_counterAddrOne[10:0];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_4_HOLD : begin
      end
      controlStateMachine_enumDef_4_PASS : begin
      end
      controlStateMachine_enumDef_4_ONCE : begin
        if(!threeInFourOutRow) begin
          if(nextRowBuffer) begin
            if(outReachRowEnd) begin
              counterAddrOne = CICC1851_counterAddrOne_1[10:0];
            end else begin
              counterAddrOne = CICC1851_counterAddrOne_3[10:0];
            end
          end
        end
      end
      controlStateMachine_enumDef_4_TWICE : begin
        if(outReachFinalRow) begin
          if(nextRowBuffer) begin
            if(!outReachRowEnd) begin
              counterAddrOne = CICC1851_counterAddrOne_5[10:0];
            end
          end
        end else begin
          if(nextRowBuffer) begin
            if(outReachRowEnd) begin
              counterAddrOne = CICC1851_counterAddrOne_9[10:0];
            end else begin
              counterAddrOne = CICC1851_counterAddrOne_11[10:0];
            end
          end else begin
            counterAddrOne = CICC1851_counterAddrOne_15[10:0];
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    mainAddrTwo = CICC1851_mainAddrTwo[10:0];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_4_HOLD : begin
      end
      controlStateMachine_enumDef_4_PASS : begin
        if(!twoInFourOutRow) begin
          if(oneInFourOutRow) begin
            if(!nextRowBuffer) begin
              if(twoInFourOutPixelAddr) begin
                mainAddrTwo = CICC1851_mainAddrTwo_1[10:0];
              end
            end
          end
        end
      end
      controlStateMachine_enumDef_4_ONCE : begin
        if(threeInFourOutRow) begin
          if(twoInFourOutPixelAddr) begin
            mainAddrTwo = CICC1851_mainAddrTwo_3[10:0];
          end
        end else begin
          if(!nextRowBuffer) begin
            mainAddrTwo = CICC1851_mainAddrTwo_5[10:0];
          end
        end
      end
      controlStateMachine_enumDef_4_TWICE : begin
        if(outReachFinalRow) begin
          if(!nextRowBuffer) begin
            if(outReachRowEnd) begin
              mainAddrTwo = CICC1851_mainAddrTwo_7[10:0];
            end else begin
              mainAddrTwo = CICC1851_mainAddrTwo_9[10:0];
            end
          end
        end else begin
          if(nextRowBuffer) begin
            if(outReachRowEnd) begin
              mainAddrTwo = CICC1851_mainAddrTwo_11[10:0];
            end else begin
              mainAddrTwo = CICC1851_mainAddrTwo_13[10:0];
            end
          end else begin
            mainAddrTwo = CICC1851_mainAddrTwo_17[10:0];
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    counterAddrTwo = CICC1851_counterAddrTwo[10:0];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_4_HOLD : begin
      end
      controlStateMachine_enumDef_4_PASS : begin
      end
      controlStateMachine_enumDef_4_ONCE : begin
        if(!threeInFourOutRow) begin
          if(!nextRowBuffer) begin
            if(outReachRowEnd) begin
              counterAddrTwo = CICC1851_counterAddrTwo_1[10:0];
            end else begin
              counterAddrTwo = CICC1851_counterAddrTwo_3[10:0];
            end
          end
        end
      end
      controlStateMachine_enumDef_4_TWICE : begin
        if(outReachFinalRow) begin
          if(!nextRowBuffer) begin
            if(!outReachRowEnd) begin
              counterAddrTwo = CICC1851_counterAddrTwo_5[10:0];
            end
          end
        end else begin
          if(nextRowBuffer) begin
            counterAddrTwo = CICC1851_counterAddrTwo_9[10:0];
          end else begin
            if(outReachRowEnd) begin
              counterAddrTwo = CICC1851_counterAddrTwo_11[10:0];
            end else begin
              counterAddrTwo = CICC1851_counterAddrTwo_13[10:0];
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign oddAddr = CICC1851_oddAddr[10:0];
  assign validStream_valid = 1'b1;
  assign CICC1851_controls_frameStart = 32'h0;
  always @(*) begin
    controls_frameStart = CICC1851_controls_frameStart[0];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_4_HOLD : begin
      end
      controlStateMachine_enumDef_4_PASS : begin
        if(frameStart) begin
          controls_frameStart = 1'b1;
        end
      end
      controlStateMachine_enumDef_4_ONCE : begin
      end
      controlStateMachine_enumDef_4_TWICE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_rowEnd = CICC1851_controls_frameStart[1];
    if(when_SuperResolutionPart2_l761) begin
      if(outReachRowEnd) begin
        controls_rowEnd = 1'b1;
      end
    end
  end

  always @(*) begin
    controls_passMode = CICC1851_controls_frameStart[2];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_4_HOLD : begin
      end
      controlStateMachine_enumDef_4_PASS : begin
        if(twoInFourOutRow) begin
          if(!when_SuperResolutionPart2_l609) begin
            if(nextRowBuffer) begin
              controls_passMode = 1'b0;
            end else begin
              controls_passMode = 1'b1;
            end
          end
        end else begin
          if(oneInFourOutRow) begin
            if(nextRowBuffer) begin
              controls_passMode = 1'b0;
            end else begin
              controls_passMode = 1'b1;
            end
          end else begin
            if(nextRowBuffer) begin
              controls_passMode = 1'b0;
            end else begin
              controls_passMode = 1'b1;
            end
          end
        end
      end
      controlStateMachine_enumDef_4_ONCE : begin
      end
      controlStateMachine_enumDef_4_TWICE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_passValid = CICC1851_controls_frameStart[3];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_4_HOLD : begin
      end
      controlStateMachine_enumDef_4_PASS : begin
        if(twoInFourOutRow) begin
          if(!when_SuperResolutionPart2_l609) begin
            controls_passValid = 1'b1;
          end
        end else begin
          if(oneInFourOutRow) begin
            controls_passValid = 1'b1;
          end else begin
            controls_passValid = 1'b1;
          end
        end
      end
      controlStateMachine_enumDef_4_ONCE : begin
      end
      controlStateMachine_enumDef_4_TWICE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_onceMode = CICC1851_controls_frameStart[6 : 4];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_4_HOLD : begin
      end
      controlStateMachine_enumDef_4_PASS : begin
      end
      controlStateMachine_enumDef_4_ONCE : begin
        if(threeInFourOutRow) begin
          if(outReachFinalRow) begin
            if(nextRowBuffer) begin
              controls_onceMode = 3'b100;
            end else begin
              controls_onceMode = 3'b101;
            end
          end else begin
            if(nextRowBuffer) begin
              controls_onceMode = {1'd0, CICC1851_controls_onceMode};
            end else begin
              controls_onceMode = {1'd0, CICC1851_controls_onceMode_1};
            end
          end
        end else begin
          if(nextRowBuffer) begin
            controls_onceMode = 3'b000;
          end else begin
            controls_onceMode = {2'd0, CICC1851_controls_onceMode_2};
          end
        end
      end
      controlStateMachine_enumDef_4_TWICE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_onceValid = CICC1851_controls_frameStart[7];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_4_HOLD : begin
      end
      controlStateMachine_enumDef_4_PASS : begin
      end
      controlStateMachine_enumDef_4_ONCE : begin
        controls_onceValid = 1'b1;
      end
      controlStateMachine_enumDef_4_TWICE : begin
      end
      default : begin
      end
    endcase
  end

  assign controls_mainCompare = CICC1851_controls_frameStart[8];
  assign controls_counterCompare = CICC1851_controls_frameStart[9];
  assign controls_mainDiff = CICC1851_controls_frameStart[17 : 10];
  assign controls_counterDiff = CICC1851_controls_frameStart[25 : 18];
  always @(*) begin
    controls_twiceCompValid = CICC1851_controls_frameStart[26];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_4_HOLD : begin
      end
      controlStateMachine_enumDef_4_PASS : begin
      end
      controlStateMachine_enumDef_4_ONCE : begin
      end
      controlStateMachine_enumDef_4_TWICE : begin
        controls_twiceCompValid = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_twiceMode = CICC1851_controls_frameStart[29 : 27];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_4_HOLD : begin
      end
      controlStateMachine_enumDef_4_PASS : begin
      end
      controlStateMachine_enumDef_4_ONCE : begin
      end
      controlStateMachine_enumDef_4_TWICE : begin
        if(outReachFinalRow) begin
          if(nextRowBuffer) begin
            if(outReachRowEnd) begin
              controls_twiceMode = 3'b100;
            end else begin
              controls_twiceMode = 3'b101;
            end
          end else begin
            if(outReachRowEnd) begin
              controls_twiceMode = {1'd0, CICC1851_controls_twiceMode};
            end else begin
              controls_twiceMode = {1'd0, CICC1851_controls_twiceMode_1};
            end
          end
        end else begin
          if(nextRowBuffer) begin
            controls_twiceMode = 3'b000;
          end else begin
            controls_twiceMode = {2'd0, CICC1851_controls_twiceMode_2};
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_inpValidFlag = CICC1851_controls_frameStart[30];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_4_HOLD : begin
        controls_inpValidFlag = 1'b1;
      end
      controlStateMachine_enumDef_4_PASS : begin
        controls_inpValidFlag = 1'b1;
      end
      controlStateMachine_enumDef_4_ONCE : begin
        controls_inpValidFlag = 1'b1;
      end
      controlStateMachine_enumDef_4_TWICE : begin
        controls_inpValidFlag = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_oddValid = CICC1851_controls_frameStart[31];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_4_HOLD : begin
      end
      controlStateMachine_enumDef_4_PASS : begin
        if(twoInFourOutRow) begin
          if(when_SuperResolutionPart2_l609) begin
            controls_oddValid = 1'b1;
          end
        end
      end
      controlStateMachine_enumDef_4_ONCE : begin
      end
      controlStateMachine_enumDef_4_TWICE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    validStream_ready = (controlStream_ready && startRead);
    validStream_ready = (mainAddrOneStream_ready && startRead);
    validStream_ready = (counterAddrOneStream_ready && startRead);
    validStream_ready = (mainAddrTwoStream_ready && startRead);
    validStream_ready = (counterAddrTwoStream_ready && startRead);
    validStream_ready = (oddAddrStream_ready && startRead);
  end

  assign controlStream_valid = (validStream_valid && startRead);
  assign controlStream_payload_frameStart = controls_frameStart;
  assign controlStream_payload_rowEnd = controls_rowEnd;
  assign controlStream_payload_passMode = controls_passMode;
  assign controlStream_payload_passValid = controls_passValid;
  assign controlStream_payload_onceMode = controls_onceMode;
  assign controlStream_payload_onceValid = controls_onceValid;
  assign controlStream_payload_mainCompare = controls_mainCompare;
  assign controlStream_payload_counterCompare = controls_counterCompare;
  assign controlStream_payload_mainDiff = controls_mainDiff;
  assign controlStream_payload_counterDiff = controls_counterDiff;
  assign controlStream_payload_twiceCompValid = controls_twiceCompValid;
  assign controlStream_payload_twiceMode = controls_twiceMode;
  assign controlStream_payload_inpValidFlag = controls_inpValidFlag;
  assign controlStream_payload_oddValid = controls_oddValid;
  assign mainAddrOneStream_valid = (validStream_valid && startRead);
  assign mainAddrOneStream_payload = mainAddrOne;
  assign counterAddrOneStream_valid = (validStream_valid && startRead);
  assign counterAddrOneStream_payload = counterAddrOne;
  assign mainAddrTwoStream_valid = (validStream_valid && startRead);
  assign mainAddrTwoStream_payload = mainAddrTwo;
  assign counterAddrTwoStream_valid = (validStream_valid && startRead);
  assign counterAddrTwoStream_payload = counterAddrTwo;
  assign oddAddrStream_valid = (validStream_valid && startRead);
  assign oddAddrStream_payload = oddAddr;
  assign pixelsIn_s2mPipe_valid = (pixelsIn_valid || pixelsIn_rValid);
  assign pixelsIn_s2mPipe_payload_pixel = (pixelsIn_rValid ? pixelsIn_rData_pixel : pixelsIn_payload_pixel);
  assign pixelsIn_s2mPipe_payload_frameStart = (pixelsIn_rValid ? pixelsIn_rData_frameStart : pixelsIn_payload_frameStart);
  assign pixelsIn_s2mPipe_payload_rowEnd = (pixelsIn_rValid ? pixelsIn_rData_rowEnd : pixelsIn_payload_rowEnd);
  always @(*) begin
    pixelsIn_s2mPipe_ready = pixelsIn_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368) begin
      pixelsIn_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368 = (! pixelsIn_s2mPipe_m2sPipe_valid);
  assign pixelsIn_s2mPipe_m2sPipe_valid = pixelsIn_s2mPipe_rValid;
  assign pixelsIn_s2mPipe_m2sPipe_payload_pixel = pixelsIn_s2mPipe_rData_pixel;
  assign pixelsIn_s2mPipe_m2sPipe_payload_frameStart = pixelsIn_s2mPipe_rData_frameStart;
  assign pixelsIn_s2mPipe_m2sPipe_payload_rowEnd = pixelsIn_s2mPipe_rData_rowEnd;
  assign passPixels_valid = (pixelsIn_s2mPipe_m2sPipe_valid && bufferEnable);
  assign pixelsIn_s2mPipe_m2sPipe_ready = (passPixels_ready && bufferEnable);
  assign passPixels_payload_pixel = pixelsIn_s2mPipe_m2sPipe_payload_pixel;
  assign passPixels_payload_frameStart = pixelsIn_s2mPipe_m2sPipe_payload_frameStart;
  assign passPixels_payload_rowEnd = pixelsIn_s2mPipe_m2sPipe_payload_rowEnd;
  assign passPixels_ready = 1'b1;
  assign passPixels_fire = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart2_l181 = ((CICC1851_when_SuperResolutionPart2_l181 == CICC1851_when_SuperResolutionPart2_l181_1) && passPixels_fire);
  assign passPixels_fire_1 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart2_l182 = (((CICC1851_when_SuperResolutionPart2_l182 == CICC1851_when_SuperResolutionPart2_l182_1) && bufferReachRowEnd) && passPixels_fire_1);
  assign passPixels_fire_2 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart2_l185 = (passPixels_payload_rowEnd && passPixels_fire_2);
  assign when_SuperResolutionPart2_l195 = (CICC1851_when_SuperResolutionPart2_l195 == 11'h0);
  assign passPixels_fire_3 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart2_l200 = (passPixels_payload_rowEnd && passPixels_fire_3);
  assign when_SuperResolutionPart2_l201 = ((bufferSwitch == 2'b10) || (bufferSwitch == 2'b00));
  assign passPixels_fire_4 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart2_l207 = (((bufferRowCount_value != 11'h0) && passPixels_payload_rowEnd) && passPixels_fire_4);
  assign when_SuperResolutionPart2_l208 = (bufferSwitch != 2'b01);
  assign when_SuperResolutionPart2_l212 = (bufferReachFinalRow && bufferReachRowEnd);
  assign controlStream_fire = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart2_l218 = (((CICC1851_when_SuperResolutionPart2_l218 == 12'h003) && controlStream_payload_rowEnd) && controlStream_fire);
  assign when_SuperResolutionPart2_l220 = 1'b1;
  assign passPixels_fire_5 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart2_l224 = (passPixels_payload_frameStart && passPixels_fire_5);
  assign pixelsOut_fire = (pixelsOut_valid && pixelsOut_ready);
  assign when_SuperResolutionPart2_l234 = ((CICC1851_when_SuperResolutionPart2_l234 == CICC1851_when_SuperResolutionPart2_l234_1) && pixelsOut_fire);
  assign pixelsOut_fire_1 = (pixelsOut_valid && pixelsOut_ready);
  assign when_SuperResolutionPart2_l235 = (((CICC1851_when_SuperResolutionPart2_l235 == CICC1851_when_SuperResolutionPart2_l235_1) && alreadyReachRowEnd) && pixelsOut_fire_1);
  assign pixelsOut_fire_2 = (pixelsOut_valid && pixelsOut_ready);
  assign pixelsOut_fire_3 = (pixelsOut_valid && pixelsOut_ready);
  assign when_SuperResolutionPart2_l246 = ((alreadyReachFinalRow && alreadyReachRowEnd) && pixelsOut_fire_3);
  assign passPixels_fire_6 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_7 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_8 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_9 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_10 = (passPixels_valid && passPixels_ready);
  assign controlStream_fire_1 = (controlStream_valid && controlStream_ready);
  assign pushing = (passPixels_fire_10 && (! controlStream_fire_1));
  assign passPixels_fire_11 = (passPixels_valid && passPixels_ready);
  assign controlStream_fire_2 = (controlStream_valid && controlStream_ready);
  assign poping = ((! passPixels_fire_11) && controlStream_fire_2);
  assign passPixels_fire_12 = (passPixels_valid && passPixels_ready);
  assign controlStream_fire_3 = (controlStream_valid && controlStream_ready);
  assign pushAndPoping = (passPixels_fire_12 && controlStream_fire_3);
  assign mainAddrOneStream_ready = (! mainAddrOneStream_rValid);
  assign mainAddrOneStream_s2mPipe_valid = (mainAddrOneStream_valid || mainAddrOneStream_rValid);
  assign mainAddrOneStream_s2mPipe_payload = (mainAddrOneStream_rValid ? mainAddrOneStream_rData : mainAddrOneStream_payload);
  always @(*) begin
    mainAddrOneStream_s2mPipe_ready = mainAddrOneStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_1) begin
      mainAddrOneStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_1 = (! mainAddrOneStream_s2mPipe_m2sPipe_valid);
  assign mainAddrOneStream_s2mPipe_m2sPipe_valid = mainAddrOneStream_s2mPipe_rValid;
  assign mainAddrOneStream_s2mPipe_m2sPipe_payload = mainAddrOneStream_s2mPipe_rData;
  assign mainAddrOneStream_s2mPipe_m2sPipe_ready = ((! CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready) || CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready = CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_mainOnePixelStream_payload = CICC1851_lineBufferOne_port1;
  assign CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_1 = readStage_mainOnePixelStream_ready;
    if(when_Stream_l368_2) begin
      CICC1851_1 = 1'b1;
    end
  end

  assign when_Stream_l368_2 = (! readStage_mainOnePixelStream_valid);
  assign readStage_mainOnePixelStream_valid = CICC1851_readStage_mainOnePixelStream_valid;
  assign readStage_mainOnePixelStream_payload = CICC1851_readStage_mainOnePixelStream_payload_2;
  assign counterAddrOneStream_ready = (! counterAddrOneStream_rValid);
  assign counterAddrOneStream_s2mPipe_valid = (counterAddrOneStream_valid || counterAddrOneStream_rValid);
  assign counterAddrOneStream_s2mPipe_payload = (counterAddrOneStream_rValid ? counterAddrOneStream_rData : counterAddrOneStream_payload);
  always @(*) begin
    counterAddrOneStream_s2mPipe_ready = counterAddrOneStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_3) begin
      counterAddrOneStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_3 = (! counterAddrOneStream_s2mPipe_m2sPipe_valid);
  assign counterAddrOneStream_s2mPipe_m2sPipe_valid = counterAddrOneStream_s2mPipe_rValid;
  assign counterAddrOneStream_s2mPipe_m2sPipe_payload = counterAddrOneStream_s2mPipe_rData;
  assign counterAddrOneStream_s2mPipe_m2sPipe_ready = ((! CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready) || CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready = CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_counterOnePixelStream_payload = CICC1851_lineBufferOne_port2;
  assign CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_2 = readStage_counterOnePixelStream_ready;
    if(when_Stream_l368_4) begin
      CICC1851_2 = 1'b1;
    end
  end

  assign when_Stream_l368_4 = (! readStage_counterOnePixelStream_valid);
  assign readStage_counterOnePixelStream_valid = CICC1851_readStage_counterOnePixelStream_valid;
  assign readStage_counterOnePixelStream_payload = CICC1851_readStage_counterOnePixelStream_payload_2;
  assign mainAddrTwoStream_ready = (! mainAddrTwoStream_rValid);
  assign mainAddrTwoStream_s2mPipe_valid = (mainAddrTwoStream_valid || mainAddrTwoStream_rValid);
  assign mainAddrTwoStream_s2mPipe_payload = (mainAddrTwoStream_rValid ? mainAddrTwoStream_rData : mainAddrTwoStream_payload);
  always @(*) begin
    mainAddrTwoStream_s2mPipe_ready = mainAddrTwoStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_5) begin
      mainAddrTwoStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_5 = (! mainAddrTwoStream_s2mPipe_m2sPipe_valid);
  assign mainAddrTwoStream_s2mPipe_m2sPipe_valid = mainAddrTwoStream_s2mPipe_rValid;
  assign mainAddrTwoStream_s2mPipe_m2sPipe_payload = mainAddrTwoStream_s2mPipe_rData;
  assign mainAddrTwoStream_s2mPipe_m2sPipe_ready = ((! CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready) || CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready = CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_mainTwoPixelStream_payload = CICC1851_lineBufferTwo_port1;
  assign CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_3 = readStage_mainTwoPixelStream_ready;
    if(when_Stream_l368_6) begin
      CICC1851_3 = 1'b1;
    end
  end

  assign when_Stream_l368_6 = (! readStage_mainTwoPixelStream_valid);
  assign readStage_mainTwoPixelStream_valid = CICC1851_readStage_mainTwoPixelStream_valid;
  assign readStage_mainTwoPixelStream_payload = CICC1851_readStage_mainTwoPixelStream_payload_2;
  assign counterAddrTwoStream_ready = (! counterAddrTwoStream_rValid);
  assign counterAddrTwoStream_s2mPipe_valid = (counterAddrTwoStream_valid || counterAddrTwoStream_rValid);
  assign counterAddrTwoStream_s2mPipe_payload = (counterAddrTwoStream_rValid ? counterAddrTwoStream_rData : counterAddrTwoStream_payload);
  always @(*) begin
    counterAddrTwoStream_s2mPipe_ready = counterAddrTwoStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_7) begin
      counterAddrTwoStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_7 = (! counterAddrTwoStream_s2mPipe_m2sPipe_valid);
  assign counterAddrTwoStream_s2mPipe_m2sPipe_valid = counterAddrTwoStream_s2mPipe_rValid;
  assign counterAddrTwoStream_s2mPipe_m2sPipe_payload = counterAddrTwoStream_s2mPipe_rData;
  assign counterAddrTwoStream_s2mPipe_m2sPipe_ready = ((! CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready) || CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready = CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_counterTwoPixelStream_payload = CICC1851_lineBufferTwo_port2;
  assign CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_4 = readStage_counterTwoPixelStream_ready;
    if(when_Stream_l368_8) begin
      CICC1851_4 = 1'b1;
    end
  end

  assign when_Stream_l368_8 = (! readStage_counterTwoPixelStream_valid);
  assign readStage_counterTwoPixelStream_valid = CICC1851_readStage_counterTwoPixelStream_valid;
  assign readStage_counterTwoPixelStream_payload = CICC1851_readStage_counterTwoPixelStream_payload_2;
  assign oddAddrStream_ready = (! oddAddrStream_rValid);
  assign oddAddrStream_s2mPipe_valid = (oddAddrStream_valid || oddAddrStream_rValid);
  assign oddAddrStream_s2mPipe_payload = (oddAddrStream_rValid ? oddAddrStream_rData : oddAddrStream_payload);
  always @(*) begin
    oddAddrStream_s2mPipe_ready = oddAddrStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_9) begin
      oddAddrStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_9 = (! oddAddrStream_s2mPipe_m2sPipe_valid);
  assign oddAddrStream_s2mPipe_m2sPipe_valid = oddAddrStream_s2mPipe_rValid;
  assign oddAddrStream_s2mPipe_m2sPipe_payload = oddAddrStream_s2mPipe_rData;
  assign oddAddrStream_s2mPipe_m2sPipe_ready = ((! CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready) || CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready = CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_oddRowPixelStream_payload = CICC1851_lineBufferOdd_port1;
  assign CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_5 = readStage_oddRowPixelStream_ready;
    if(when_Stream_l368_10) begin
      CICC1851_5 = 1'b1;
    end
  end

  assign when_Stream_l368_10 = (! readStage_oddRowPixelStream_valid);
  assign readStage_oddRowPixelStream_valid = CICC1851_readStage_oddRowPixelStream_valid;
  assign readStage_oddRowPixelStream_payload = CICC1851_readStage_oddRowPixelStream_payload_2;
  assign controlStream_ready = (! controlStream_rValid);
  assign controlStream_s2mPipe_valid = (controlStream_valid || controlStream_rValid);
  assign controlStream_s2mPipe_payload_frameStart = (controlStream_rValid ? controlStream_rData_frameStart : controlStream_payload_frameStart);
  assign controlStream_s2mPipe_payload_rowEnd = (controlStream_rValid ? controlStream_rData_rowEnd : controlStream_payload_rowEnd);
  assign controlStream_s2mPipe_payload_passMode = (controlStream_rValid ? controlStream_rData_passMode : controlStream_payload_passMode);
  assign controlStream_s2mPipe_payload_passValid = (controlStream_rValid ? controlStream_rData_passValid : controlStream_payload_passValid);
  assign controlStream_s2mPipe_payload_onceMode = (controlStream_rValid ? controlStream_rData_onceMode : controlStream_payload_onceMode);
  assign controlStream_s2mPipe_payload_onceValid = (controlStream_rValid ? controlStream_rData_onceValid : controlStream_payload_onceValid);
  assign controlStream_s2mPipe_payload_mainCompare = (controlStream_rValid ? controlStream_rData_mainCompare : controlStream_payload_mainCompare);
  assign controlStream_s2mPipe_payload_counterCompare = (controlStream_rValid ? controlStream_rData_counterCompare : controlStream_payload_counterCompare);
  assign controlStream_s2mPipe_payload_mainDiff = (controlStream_rValid ? controlStream_rData_mainDiff : controlStream_payload_mainDiff);
  assign controlStream_s2mPipe_payload_counterDiff = (controlStream_rValid ? controlStream_rData_counterDiff : controlStream_payload_counterDiff);
  assign controlStream_s2mPipe_payload_twiceCompValid = (controlStream_rValid ? controlStream_rData_twiceCompValid : controlStream_payload_twiceCompValid);
  assign controlStream_s2mPipe_payload_twiceMode = (controlStream_rValid ? controlStream_rData_twiceMode : controlStream_payload_twiceMode);
  assign controlStream_s2mPipe_payload_inpValidFlag = (controlStream_rValid ? controlStream_rData_inpValidFlag : controlStream_payload_inpValidFlag);
  assign controlStream_s2mPipe_payload_oddValid = (controlStream_rValid ? controlStream_rData_oddValid : controlStream_payload_oddValid);
  always @(*) begin
    controlStream_s2mPipe_ready = controlStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_11) begin
      controlStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_11 = (! controlStream_s2mPipe_m2sPipe_valid);
  assign controlStream_s2mPipe_m2sPipe_valid = controlStream_s2mPipe_rValid;
  assign controlStream_s2mPipe_m2sPipe_payload_frameStart = controlStream_s2mPipe_rData_frameStart;
  assign controlStream_s2mPipe_m2sPipe_payload_rowEnd = controlStream_s2mPipe_rData_rowEnd;
  assign controlStream_s2mPipe_m2sPipe_payload_passMode = controlStream_s2mPipe_rData_passMode;
  assign controlStream_s2mPipe_m2sPipe_payload_passValid = controlStream_s2mPipe_rData_passValid;
  assign controlStream_s2mPipe_m2sPipe_payload_onceMode = controlStream_s2mPipe_rData_onceMode;
  assign controlStream_s2mPipe_m2sPipe_payload_onceValid = controlStream_s2mPipe_rData_onceValid;
  assign controlStream_s2mPipe_m2sPipe_payload_mainCompare = controlStream_s2mPipe_rData_mainCompare;
  assign controlStream_s2mPipe_m2sPipe_payload_counterCompare = controlStream_s2mPipe_rData_counterCompare;
  assign controlStream_s2mPipe_m2sPipe_payload_mainDiff = controlStream_s2mPipe_rData_mainDiff;
  assign controlStream_s2mPipe_m2sPipe_payload_counterDiff = controlStream_s2mPipe_rData_counterDiff;
  assign controlStream_s2mPipe_m2sPipe_payload_twiceCompValid = controlStream_s2mPipe_rData_twiceCompValid;
  assign controlStream_s2mPipe_m2sPipe_payload_twiceMode = controlStream_s2mPipe_rData_twiceMode;
  assign controlStream_s2mPipe_m2sPipe_payload_inpValidFlag = controlStream_s2mPipe_rData_inpValidFlag;
  assign controlStream_s2mPipe_m2sPipe_payload_oddValid = controlStream_s2mPipe_rData_oddValid;
  always @(*) begin
    controlStream_s2mPipe_m2sPipe_ready = controlStream_s2mPipe_m2sPipe_m2sPipe_ready;
    if(when_Stream_l368_12) begin
      controlStream_s2mPipe_m2sPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_12 = (! controlStream_s2mPipe_m2sPipe_m2sPipe_valid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_valid = controlStream_s2mPipe_m2sPipe_rValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_frameStart = controlStream_s2mPipe_m2sPipe_rData_frameStart;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_rowEnd = controlStream_s2mPipe_m2sPipe_rData_rowEnd;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passMode = controlStream_s2mPipe_m2sPipe_rData_passMode;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passValid = controlStream_s2mPipe_m2sPipe_rData_passValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceMode = controlStream_s2mPipe_m2sPipe_rData_onceMode;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceValid = controlStream_s2mPipe_m2sPipe_rData_onceValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainCompare = controlStream_s2mPipe_m2sPipe_rData_mainCompare;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterCompare = controlStream_s2mPipe_m2sPipe_rData_counterCompare;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDiff = controlStream_s2mPipe_m2sPipe_rData_mainDiff;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDiff = controlStream_s2mPipe_m2sPipe_rData_counterDiff;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceCompValid = controlStream_s2mPipe_m2sPipe_rData_twiceCompValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceMode = controlStream_s2mPipe_m2sPipe_rData_twiceMode;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_inpValidFlag = controlStream_s2mPipe_m2sPipe_rData_inpValidFlag;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_oddValid = controlStream_s2mPipe_m2sPipe_rData_oddValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_ready = (! controlStream_s2mPipe_m2sPipe_m2sPipe_rValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_valid = (controlStream_s2mPipe_m2sPipe_m2sPipe_valid || controlStream_s2mPipe_m2sPipe_m2sPipe_rValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_frameStart = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_frameStart : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_frameStart);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_rowEnd = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_rowEnd : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_rowEnd);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_passMode = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_passMode : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passMode);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_passValid = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_passValid : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_onceMode = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_onceMode : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceMode);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_onceValid = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_onceValid : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainCompare = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainCompare : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainCompare);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterCompare = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterCompare : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterCompare);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainDiff = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainDiff : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDiff);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterDiff = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterDiff : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDiff);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_twiceCompValid = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_twiceCompValid : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceCompValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_twiceMode = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_twiceMode : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceMode);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_inpValidFlag = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_inpValidFlag : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_inpValidFlag);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_oddValid = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_oddValid : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_oddValid);
  always @(*) begin
    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready = readStage_controlPipe_ready;
    if(when_Stream_l368_13) begin
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_13 = (! readStage_controlPipe_valid);
  assign readStage_controlPipe_valid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rValid;
  assign readStage_controlPipe_payload_frameStart = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_frameStart;
  assign readStage_controlPipe_payload_rowEnd = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_rowEnd;
  assign readStage_controlPipe_payload_passMode = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_passMode;
  assign readStage_controlPipe_payload_passValid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_passValid;
  assign readStage_controlPipe_payload_onceMode = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_onceMode;
  assign readStage_controlPipe_payload_onceValid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_onceValid;
  assign readStage_controlPipe_payload_mainCompare = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainCompare;
  assign readStage_controlPipe_payload_counterCompare = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterCompare;
  assign readStage_controlPipe_payload_mainDiff = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainDiff;
  assign readStage_controlPipe_payload_counterDiff = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterDiff;
  assign readStage_controlPipe_payload_twiceCompValid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_twiceCompValid;
  assign readStage_controlPipe_payload_twiceMode = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_twiceMode;
  assign readStage_controlPipe_payload_inpValidFlag = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_inpValidFlag;
  assign readStage_controlPipe_payload_oddValid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_oddValid;
  assign readStage_mainOnePixelStream_ready = (! readStage_mainOnePixelStream_rValid);
  assign readStage_mainOnePixelStream_s2mPipe_valid = (readStage_mainOnePixelStream_valid || readStage_mainOnePixelStream_rValid);
  assign readStage_mainOnePixelStream_s2mPipe_payload = (readStage_mainOnePixelStream_rValid ? readStage_mainOnePixelStream_rData : readStage_mainOnePixelStream_payload);
  always @(*) begin
    readStage_mainOnePixelStream_s2mPipe_ready = compareStage_mainOnePixelStream_ready;
    if(when_Stream_l368_14) begin
      readStage_mainOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_14 = (! compareStage_mainOnePixelStream_valid);
  assign compareStage_mainOnePixelStream_valid = readStage_mainOnePixelStream_s2mPipe_rValid;
  assign compareStage_mainOnePixelStream_payload = readStage_mainOnePixelStream_s2mPipe_rData;
  assign readStage_counterOnePixelStream_ready = (! readStage_counterOnePixelStream_rValid);
  assign readStage_counterOnePixelStream_s2mPipe_valid = (readStage_counterOnePixelStream_valid || readStage_counterOnePixelStream_rValid);
  assign readStage_counterOnePixelStream_s2mPipe_payload = (readStage_counterOnePixelStream_rValid ? readStage_counterOnePixelStream_rData : readStage_counterOnePixelStream_payload);
  always @(*) begin
    readStage_counterOnePixelStream_s2mPipe_ready = compareStage_counterOnePixelStream_ready;
    if(when_Stream_l368_15) begin
      readStage_counterOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_15 = (! compareStage_counterOnePixelStream_valid);
  assign compareStage_counterOnePixelStream_valid = readStage_counterOnePixelStream_s2mPipe_rValid;
  assign compareStage_counterOnePixelStream_payload = readStage_counterOnePixelStream_s2mPipe_rData;
  assign readStage_mainTwoPixelStream_ready = (! readStage_mainTwoPixelStream_rValid);
  assign readStage_mainTwoPixelStream_s2mPipe_valid = (readStage_mainTwoPixelStream_valid || readStage_mainTwoPixelStream_rValid);
  assign readStage_mainTwoPixelStream_s2mPipe_payload = (readStage_mainTwoPixelStream_rValid ? readStage_mainTwoPixelStream_rData : readStage_mainTwoPixelStream_payload);
  always @(*) begin
    readStage_mainTwoPixelStream_s2mPipe_ready = compareStage_mainTwoPixelStream_ready;
    if(when_Stream_l368_16) begin
      readStage_mainTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_16 = (! compareStage_mainTwoPixelStream_valid);
  assign compareStage_mainTwoPixelStream_valid = readStage_mainTwoPixelStream_s2mPipe_rValid;
  assign compareStage_mainTwoPixelStream_payload = readStage_mainTwoPixelStream_s2mPipe_rData;
  assign readStage_counterTwoPixelStream_ready = (! readStage_counterTwoPixelStream_rValid);
  assign readStage_counterTwoPixelStream_s2mPipe_valid = (readStage_counterTwoPixelStream_valid || readStage_counterTwoPixelStream_rValid);
  assign readStage_counterTwoPixelStream_s2mPipe_payload = (readStage_counterTwoPixelStream_rValid ? readStage_counterTwoPixelStream_rData : readStage_counterTwoPixelStream_payload);
  always @(*) begin
    readStage_counterTwoPixelStream_s2mPipe_ready = compareStage_counterTwoPixelStream_ready;
    if(when_Stream_l368_17) begin
      readStage_counterTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_17 = (! compareStage_counterTwoPixelStream_valid);
  assign compareStage_counterTwoPixelStream_valid = readStage_counterTwoPixelStream_s2mPipe_rValid;
  assign compareStage_counterTwoPixelStream_payload = readStage_counterTwoPixelStream_s2mPipe_rData;
  assign readStage_oddRowPixelStream_ready = (! readStage_oddRowPixelStream_rValid);
  assign readStage_oddRowPixelStream_s2mPipe_valid = (readStage_oddRowPixelStream_valid || readStage_oddRowPixelStream_rValid);
  assign readStage_oddRowPixelStream_s2mPipe_payload = (readStage_oddRowPixelStream_rValid ? readStage_oddRowPixelStream_rData : readStage_oddRowPixelStream_payload);
  always @(*) begin
    readStage_oddRowPixelStream_s2mPipe_ready = compareStage_oddRowPixelStream_ready;
    if(when_Stream_l368_18) begin
      readStage_oddRowPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_18 = (! compareStage_oddRowPixelStream_valid);
  assign compareStage_oddRowPixelStream_valid = readStage_oddRowPixelStream_s2mPipe_rValid;
  assign compareStage_oddRowPixelStream_payload = readStage_oddRowPixelStream_s2mPipe_rData;
  always @(*) begin
    CICC1851_readStage_controlPipe_translated_payload_mainCompare = readStage_controlPipe_payload_mainCompare;
    if(readStage_controlPipe_payload_onceValid) begin
      case(readStage_controlPipe_payload_onceMode)
        3'b000 : begin
          if(when_SuperResolutionPart2_l290) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        3'b001 : begin
          if(when_SuperResolutionPart2_l294) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        3'b010 : begin
          if(when_SuperResolutionPart2_l298) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        3'b011 : begin
          if(when_SuperResolutionPart2_l302) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        3'b100 : begin
          CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
        end
        3'b101 : begin
          CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
        end
        default : begin
        end
      endcase
    end
    if(readStage_controlPipe_payload_twiceCompValid) begin
      case(readStage_controlPipe_payload_twiceMode)
        3'b000 : begin
          if(when_SuperResolutionPart2_l313) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        3'b001 : begin
          if(when_SuperResolutionPart2_l319) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        3'b010 : begin
          CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
        end
        3'b011 : begin
          if(when_SuperResolutionPart2_l326) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        3'b100 : begin
          CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
        end
        3'b101 : begin
          if(when_SuperResolutionPart2_l331) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    CICC1851_readStage_controlPipe_translated_payload_counterCompare = readStage_controlPipe_payload_counterCompare;
    if(readStage_controlPipe_payload_twiceCompValid) begin
      case(readStage_controlPipe_payload_twiceMode)
        3'b000 : begin
          if(when_SuperResolutionPart2_l315) begin
            CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
          end
        end
        3'b001 : begin
          if(when_SuperResolutionPart2_l321) begin
            CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
          end
        end
        default : begin
        end
      endcase
    end
  end

  assign when_SuperResolutionPart2_l290 = (readStage_counterOnePixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart2_l294 = (readStage_counterTwoPixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart2_l298 = (readStage_mainTwoPixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart2_l302 = (readStage_mainOnePixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart2_l313 = (readStage_mainTwoPixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart2_l315 = (readStage_counterOnePixelStream_payload <= readStage_counterTwoPixelStream_payload);
  assign when_SuperResolutionPart2_l319 = (readStage_mainOnePixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart2_l321 = (readStage_counterTwoPixelStream_payload <= readStage_counterOnePixelStream_payload);
  assign when_SuperResolutionPart2_l326 = (readStage_counterTwoPixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart2_l331 = (readStage_counterOnePixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign readStage_controlPipe_translated_valid = readStage_controlPipe_valid;
  assign readStage_controlPipe_ready = readStage_controlPipe_translated_ready;
  assign readStage_controlPipe_translated_payload_frameStart = readStage_controlPipe_payload_frameStart;
  assign readStage_controlPipe_translated_payload_rowEnd = readStage_controlPipe_payload_rowEnd;
  assign readStage_controlPipe_translated_payload_passMode = readStage_controlPipe_payload_passMode;
  assign readStage_controlPipe_translated_payload_passValid = readStage_controlPipe_payload_passValid;
  assign readStage_controlPipe_translated_payload_onceMode = readStage_controlPipe_payload_onceMode;
  assign readStage_controlPipe_translated_payload_onceValid = readStage_controlPipe_payload_onceValid;
  assign readStage_controlPipe_translated_payload_mainCompare = CICC1851_readStage_controlPipe_translated_payload_mainCompare;
  assign readStage_controlPipe_translated_payload_counterCompare = CICC1851_readStage_controlPipe_translated_payload_counterCompare;
  assign readStage_controlPipe_translated_payload_mainDiff = readStage_controlPipe_payload_mainDiff;
  assign readStage_controlPipe_translated_payload_counterDiff = readStage_controlPipe_payload_counterDiff;
  assign readStage_controlPipe_translated_payload_twiceCompValid = readStage_controlPipe_payload_twiceCompValid;
  assign readStage_controlPipe_translated_payload_twiceMode = readStage_controlPipe_payload_twiceMode;
  assign readStage_controlPipe_translated_payload_inpValidFlag = readStage_controlPipe_payload_inpValidFlag;
  assign readStage_controlPipe_translated_payload_oddValid = readStage_controlPipe_payload_oddValid;
  assign readStage_controlPipe_translated_ready = (! readStage_controlPipe_translated_rValid);
  assign readStage_controlPipe_translated_s2mPipe_valid = (readStage_controlPipe_translated_valid || readStage_controlPipe_translated_rValid);
  assign readStage_controlPipe_translated_s2mPipe_payload_frameStart = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_frameStart : readStage_controlPipe_translated_payload_frameStart);
  assign readStage_controlPipe_translated_s2mPipe_payload_rowEnd = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_rowEnd : readStage_controlPipe_translated_payload_rowEnd);
  assign readStage_controlPipe_translated_s2mPipe_payload_passMode = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_passMode : readStage_controlPipe_translated_payload_passMode);
  assign readStage_controlPipe_translated_s2mPipe_payload_passValid = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_passValid : readStage_controlPipe_translated_payload_passValid);
  assign readStage_controlPipe_translated_s2mPipe_payload_onceMode = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_onceMode : readStage_controlPipe_translated_payload_onceMode);
  assign readStage_controlPipe_translated_s2mPipe_payload_onceValid = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_onceValid : readStage_controlPipe_translated_payload_onceValid);
  assign readStage_controlPipe_translated_s2mPipe_payload_mainCompare = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_mainCompare : readStage_controlPipe_translated_payload_mainCompare);
  assign readStage_controlPipe_translated_s2mPipe_payload_counterCompare = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_counterCompare : readStage_controlPipe_translated_payload_counterCompare);
  assign readStage_controlPipe_translated_s2mPipe_payload_mainDiff = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_mainDiff : readStage_controlPipe_translated_payload_mainDiff);
  assign readStage_controlPipe_translated_s2mPipe_payload_counterDiff = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_counterDiff : readStage_controlPipe_translated_payload_counterDiff);
  assign readStage_controlPipe_translated_s2mPipe_payload_twiceCompValid = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_twiceCompValid : readStage_controlPipe_translated_payload_twiceCompValid);
  assign readStage_controlPipe_translated_s2mPipe_payload_twiceMode = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_twiceMode : readStage_controlPipe_translated_payload_twiceMode);
  assign readStage_controlPipe_translated_s2mPipe_payload_inpValidFlag = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_inpValidFlag : readStage_controlPipe_translated_payload_inpValidFlag);
  assign readStage_controlPipe_translated_s2mPipe_payload_oddValid = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_oddValid : readStage_controlPipe_translated_payload_oddValid);
  always @(*) begin
    readStage_controlPipe_translated_s2mPipe_ready = compareStage_controlPipe_ready;
    if(when_Stream_l368_19) begin
      readStage_controlPipe_translated_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_19 = (! compareStage_controlPipe_valid);
  assign compareStage_controlPipe_valid = readStage_controlPipe_translated_s2mPipe_rValid;
  assign compareStage_controlPipe_payload_frameStart = readStage_controlPipe_translated_s2mPipe_rData_frameStart;
  assign compareStage_controlPipe_payload_rowEnd = readStage_controlPipe_translated_s2mPipe_rData_rowEnd;
  assign compareStage_controlPipe_payload_passMode = readStage_controlPipe_translated_s2mPipe_rData_passMode;
  assign compareStage_controlPipe_payload_passValid = readStage_controlPipe_translated_s2mPipe_rData_passValid;
  assign compareStage_controlPipe_payload_onceMode = readStage_controlPipe_translated_s2mPipe_rData_onceMode;
  assign compareStage_controlPipe_payload_onceValid = readStage_controlPipe_translated_s2mPipe_rData_onceValid;
  assign compareStage_controlPipe_payload_mainCompare = readStage_controlPipe_translated_s2mPipe_rData_mainCompare;
  assign compareStage_controlPipe_payload_counterCompare = readStage_controlPipe_translated_s2mPipe_rData_counterCompare;
  assign compareStage_controlPipe_payload_mainDiff = readStage_controlPipe_translated_s2mPipe_rData_mainDiff;
  assign compareStage_controlPipe_payload_counterDiff = readStage_controlPipe_translated_s2mPipe_rData_counterDiff;
  assign compareStage_controlPipe_payload_twiceCompValid = readStage_controlPipe_translated_s2mPipe_rData_twiceCompValid;
  assign compareStage_controlPipe_payload_twiceMode = readStage_controlPipe_translated_s2mPipe_rData_twiceMode;
  assign compareStage_controlPipe_payload_inpValidFlag = readStage_controlPipe_translated_s2mPipe_rData_inpValidFlag;
  assign compareStage_controlPipe_payload_oddValid = readStage_controlPipe_translated_s2mPipe_rData_oddValid;
  assign compareStage_mainOnePixelStream_ready = (! compareStage_mainOnePixelStream_rValid);
  assign compareStage_mainOnePixelStream_s2mPipe_valid = (compareStage_mainOnePixelStream_valid || compareStage_mainOnePixelStream_rValid);
  assign compareStage_mainOnePixelStream_s2mPipe_payload = (compareStage_mainOnePixelStream_rValid ? compareStage_mainOnePixelStream_rData : compareStage_mainOnePixelStream_payload);
  always @(*) begin
    compareStage_mainOnePixelStream_s2mPipe_ready = diffStage_mainOnePixelStream_ready;
    if(when_Stream_l368_20) begin
      compareStage_mainOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_20 = (! diffStage_mainOnePixelStream_valid);
  assign diffStage_mainOnePixelStream_valid = compareStage_mainOnePixelStream_s2mPipe_rValid;
  assign diffStage_mainOnePixelStream_payload = compareStage_mainOnePixelStream_s2mPipe_rData;
  assign compareStage_counterOnePixelStream_ready = (! compareStage_counterOnePixelStream_rValid);
  assign compareStage_counterOnePixelStream_s2mPipe_valid = (compareStage_counterOnePixelStream_valid || compareStage_counterOnePixelStream_rValid);
  assign compareStage_counterOnePixelStream_s2mPipe_payload = (compareStage_counterOnePixelStream_rValid ? compareStage_counterOnePixelStream_rData : compareStage_counterOnePixelStream_payload);
  always @(*) begin
    compareStage_counterOnePixelStream_s2mPipe_ready = diffStage_counterOnePixelStream_ready;
    if(when_Stream_l368_21) begin
      compareStage_counterOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_21 = (! diffStage_counterOnePixelStream_valid);
  assign diffStage_counterOnePixelStream_valid = compareStage_counterOnePixelStream_s2mPipe_rValid;
  assign diffStage_counterOnePixelStream_payload = compareStage_counterOnePixelStream_s2mPipe_rData;
  assign compareStage_mainTwoPixelStream_ready = (! compareStage_mainTwoPixelStream_rValid);
  assign compareStage_mainTwoPixelStream_s2mPipe_valid = (compareStage_mainTwoPixelStream_valid || compareStage_mainTwoPixelStream_rValid);
  assign compareStage_mainTwoPixelStream_s2mPipe_payload = (compareStage_mainTwoPixelStream_rValid ? compareStage_mainTwoPixelStream_rData : compareStage_mainTwoPixelStream_payload);
  always @(*) begin
    compareStage_mainTwoPixelStream_s2mPipe_ready = diffStage_mainTwoPixelStream_ready;
    if(when_Stream_l368_22) begin
      compareStage_mainTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_22 = (! diffStage_mainTwoPixelStream_valid);
  assign diffStage_mainTwoPixelStream_valid = compareStage_mainTwoPixelStream_s2mPipe_rValid;
  assign diffStage_mainTwoPixelStream_payload = compareStage_mainTwoPixelStream_s2mPipe_rData;
  assign compareStage_counterTwoPixelStream_ready = (! compareStage_counterTwoPixelStream_rValid);
  assign compareStage_counterTwoPixelStream_s2mPipe_valid = (compareStage_counterTwoPixelStream_valid || compareStage_counterTwoPixelStream_rValid);
  assign compareStage_counterTwoPixelStream_s2mPipe_payload = (compareStage_counterTwoPixelStream_rValid ? compareStage_counterTwoPixelStream_rData : compareStage_counterTwoPixelStream_payload);
  always @(*) begin
    compareStage_counterTwoPixelStream_s2mPipe_ready = diffStage_counterTwoPixelStream_ready;
    if(when_Stream_l368_23) begin
      compareStage_counterTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_23 = (! diffStage_counterTwoPixelStream_valid);
  assign diffStage_counterTwoPixelStream_valid = compareStage_counterTwoPixelStream_s2mPipe_rValid;
  assign diffStage_counterTwoPixelStream_payload = compareStage_counterTwoPixelStream_s2mPipe_rData;
  assign compareStage_oddRowPixelStream_ready = (! compareStage_oddRowPixelStream_rValid);
  assign compareStage_oddRowPixelStream_s2mPipe_valid = (compareStage_oddRowPixelStream_valid || compareStage_oddRowPixelStream_rValid);
  assign compareStage_oddRowPixelStream_s2mPipe_payload = (compareStage_oddRowPixelStream_rValid ? compareStage_oddRowPixelStream_rData : compareStage_oddRowPixelStream_payload);
  always @(*) begin
    compareStage_oddRowPixelStream_s2mPipe_ready = diffStage_oddRowPixelStream_ready;
    if(when_Stream_l368_24) begin
      compareStage_oddRowPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_24 = (! diffStage_oddRowPixelStream_valid);
  assign diffStage_oddRowPixelStream_valid = compareStage_oddRowPixelStream_s2mPipe_rValid;
  assign diffStage_oddRowPixelStream_payload = compareStage_oddRowPixelStream_s2mPipe_rData;
  always @(*) begin
    CICC1851_compareStage_controlPipe_translated_payload_mainDiff = compareStage_controlPipe_payload_mainDiff;
    if(compareStage_controlPipe_payload_onceValid) begin
      case(compareStage_controlPipe_payload_onceMode)
        3'b000 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_counterOnePixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterOnePixelStream_payload - compareStage_mainOnePixelStream_payload);
          end
        end
        3'b001 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterTwoPixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainTwoPixelStream_payload);
          end
        end
        3'b010 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_mainTwoPixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_mainOnePixelStream_payload);
          end
        end
        3'b011 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_mainOnePixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_mainTwoPixelStream_payload);
          end
        end
        3'b100 : begin
          CICC1851_compareStage_controlPipe_translated_payload_mainDiff = 8'h0;
        end
        3'b101 : begin
          CICC1851_compareStage_controlPipe_translated_payload_mainDiff = 8'h0;
        end
        default : begin
        end
      endcase
    end
    if(compareStage_controlPipe_payload_twiceCompValid) begin
      case(compareStage_controlPipe_payload_twiceMode)
        3'b000 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_mainTwoPixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_mainOnePixelStream_payload);
          end
        end
        3'b001 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_mainOnePixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_mainTwoPixelStream_payload);
          end
        end
        3'b010 : begin
          CICC1851_compareStage_controlPipe_translated_payload_mainDiff = 8'h0;
        end
        3'b011 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterTwoPixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainTwoPixelStream_payload);
          end
        end
        3'b100 : begin
          CICC1851_compareStage_controlPipe_translated_payload_mainDiff = 8'h0;
        end
        3'b101 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_counterOnePixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterOnePixelStream_payload - compareStage_mainOnePixelStream_payload);
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    CICC1851_compareStage_controlPipe_translated_payload_counterDiff = compareStage_controlPipe_payload_counterDiff;
    if(compareStage_controlPipe_payload_twiceCompValid) begin
      case(compareStage_controlPipe_payload_twiceMode)
        3'b000 : begin
          if(compareStage_controlPipe_payload_counterCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterTwoPixelStream_payload - compareStage_counterOnePixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterOnePixelStream_payload - compareStage_counterTwoPixelStream_payload);
          end
        end
        3'b001 : begin
          if(compareStage_controlPipe_payload_counterCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterOnePixelStream_payload - compareStage_counterTwoPixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterTwoPixelStream_payload - compareStage_counterOnePixelStream_payload);
          end
        end
        default : begin
        end
      endcase
    end
  end

  assign compareStage_controlPipe_translated_valid = compareStage_controlPipe_valid;
  assign compareStage_controlPipe_ready = compareStage_controlPipe_translated_ready;
  assign compareStage_controlPipe_translated_payload_frameStart = compareStage_controlPipe_payload_frameStart;
  assign compareStage_controlPipe_translated_payload_rowEnd = compareStage_controlPipe_payload_rowEnd;
  assign compareStage_controlPipe_translated_payload_passMode = compareStage_controlPipe_payload_passMode;
  assign compareStage_controlPipe_translated_payload_passValid = compareStage_controlPipe_payload_passValid;
  assign compareStage_controlPipe_translated_payload_onceMode = compareStage_controlPipe_payload_onceMode;
  assign compareStage_controlPipe_translated_payload_onceValid = compareStage_controlPipe_payload_onceValid;
  assign compareStage_controlPipe_translated_payload_mainCompare = compareStage_controlPipe_payload_mainCompare;
  assign compareStage_controlPipe_translated_payload_counterCompare = compareStage_controlPipe_payload_counterCompare;
  assign compareStage_controlPipe_translated_payload_mainDiff = CICC1851_compareStage_controlPipe_translated_payload_mainDiff;
  assign compareStage_controlPipe_translated_payload_counterDiff = CICC1851_compareStage_controlPipe_translated_payload_counterDiff;
  assign compareStage_controlPipe_translated_payload_twiceCompValid = compareStage_controlPipe_payload_twiceCompValid;
  assign compareStage_controlPipe_translated_payload_twiceMode = compareStage_controlPipe_payload_twiceMode;
  assign compareStage_controlPipe_translated_payload_inpValidFlag = compareStage_controlPipe_payload_inpValidFlag;
  assign compareStage_controlPipe_translated_payload_oddValid = compareStage_controlPipe_payload_oddValid;
  assign compareStage_controlPipe_translated_ready = (! compareStage_controlPipe_translated_rValid);
  assign compareStage_controlPipe_translated_s2mPipe_valid = (compareStage_controlPipe_translated_valid || compareStage_controlPipe_translated_rValid);
  assign compareStage_controlPipe_translated_s2mPipe_payload_frameStart = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_frameStart : compareStage_controlPipe_translated_payload_frameStart);
  assign compareStage_controlPipe_translated_s2mPipe_payload_rowEnd = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_rowEnd : compareStage_controlPipe_translated_payload_rowEnd);
  assign compareStage_controlPipe_translated_s2mPipe_payload_passMode = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_passMode : compareStage_controlPipe_translated_payload_passMode);
  assign compareStage_controlPipe_translated_s2mPipe_payload_passValid = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_passValid : compareStage_controlPipe_translated_payload_passValid);
  assign compareStage_controlPipe_translated_s2mPipe_payload_onceMode = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_onceMode : compareStage_controlPipe_translated_payload_onceMode);
  assign compareStage_controlPipe_translated_s2mPipe_payload_onceValid = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_onceValid : compareStage_controlPipe_translated_payload_onceValid);
  assign compareStage_controlPipe_translated_s2mPipe_payload_mainCompare = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_mainCompare : compareStage_controlPipe_translated_payload_mainCompare);
  assign compareStage_controlPipe_translated_s2mPipe_payload_counterCompare = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_counterCompare : compareStage_controlPipe_translated_payload_counterCompare);
  assign compareStage_controlPipe_translated_s2mPipe_payload_mainDiff = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_mainDiff : compareStage_controlPipe_translated_payload_mainDiff);
  assign compareStage_controlPipe_translated_s2mPipe_payload_counterDiff = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_counterDiff : compareStage_controlPipe_translated_payload_counterDiff);
  assign compareStage_controlPipe_translated_s2mPipe_payload_twiceCompValid = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_twiceCompValid : compareStage_controlPipe_translated_payload_twiceCompValid);
  assign compareStage_controlPipe_translated_s2mPipe_payload_twiceMode = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_twiceMode : compareStage_controlPipe_translated_payload_twiceMode);
  assign compareStage_controlPipe_translated_s2mPipe_payload_inpValidFlag = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_inpValidFlag : compareStage_controlPipe_translated_payload_inpValidFlag);
  assign compareStage_controlPipe_translated_s2mPipe_payload_oddValid = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_oddValid : compareStage_controlPipe_translated_payload_oddValid);
  always @(*) begin
    compareStage_controlPipe_translated_s2mPipe_ready = diffStage_controlPipe_ready;
    if(when_Stream_l368_25) begin
      compareStage_controlPipe_translated_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_25 = (! diffStage_controlPipe_valid);
  assign diffStage_controlPipe_valid = compareStage_controlPipe_translated_s2mPipe_rValid;
  assign diffStage_controlPipe_payload_frameStart = compareStage_controlPipe_translated_s2mPipe_rData_frameStart;
  assign diffStage_controlPipe_payload_rowEnd = compareStage_controlPipe_translated_s2mPipe_rData_rowEnd;
  assign diffStage_controlPipe_payload_passMode = compareStage_controlPipe_translated_s2mPipe_rData_passMode;
  assign diffStage_controlPipe_payload_passValid = compareStage_controlPipe_translated_s2mPipe_rData_passValid;
  assign diffStage_controlPipe_payload_onceMode = compareStage_controlPipe_translated_s2mPipe_rData_onceMode;
  assign diffStage_controlPipe_payload_onceValid = compareStage_controlPipe_translated_s2mPipe_rData_onceValid;
  assign diffStage_controlPipe_payload_mainCompare = compareStage_controlPipe_translated_s2mPipe_rData_mainCompare;
  assign diffStage_controlPipe_payload_counterCompare = compareStage_controlPipe_translated_s2mPipe_rData_counterCompare;
  assign diffStage_controlPipe_payload_mainDiff = compareStage_controlPipe_translated_s2mPipe_rData_mainDiff;
  assign diffStage_controlPipe_payload_counterDiff = compareStage_controlPipe_translated_s2mPipe_rData_counterDiff;
  assign diffStage_controlPipe_payload_twiceCompValid = compareStage_controlPipe_translated_s2mPipe_rData_twiceCompValid;
  assign diffStage_controlPipe_payload_twiceMode = compareStage_controlPipe_translated_s2mPipe_rData_twiceMode;
  assign diffStage_controlPipe_payload_inpValidFlag = compareStage_controlPipe_translated_s2mPipe_rData_inpValidFlag;
  assign diffStage_controlPipe_payload_oddValid = compareStage_controlPipe_translated_s2mPipe_rData_oddValid;
  assign diffStage_mainOnePixelStream_ready = (! diffStage_mainOnePixelStream_rValid);
  assign diffStage_mainOnePixelStream_s2mPipe_valid = (diffStage_mainOnePixelStream_valid || diffStage_mainOnePixelStream_rValid);
  assign diffStage_mainOnePixelStream_s2mPipe_payload = (diffStage_mainOnePixelStream_rValid ? diffStage_mainOnePixelStream_rData : diffStage_mainOnePixelStream_payload);
  always @(*) begin
    diffStage_mainOnePixelStream_s2mPipe_ready = resultStage_mainOnePixelStream_ready;
    if(when_Stream_l368_26) begin
      diffStage_mainOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_26 = (! resultStage_mainOnePixelStream_valid);
  assign resultStage_mainOnePixelStream_valid = diffStage_mainOnePixelStream_s2mPipe_rValid;
  assign resultStage_mainOnePixelStream_payload = diffStage_mainOnePixelStream_s2mPipe_rData;
  assign diffStage_counterOnePixelStream_ready = (! diffStage_counterOnePixelStream_rValid);
  assign diffStage_counterOnePixelStream_s2mPipe_valid = (diffStage_counterOnePixelStream_valid || diffStage_counterOnePixelStream_rValid);
  assign diffStage_counterOnePixelStream_s2mPipe_payload = (diffStage_counterOnePixelStream_rValid ? diffStage_counterOnePixelStream_rData : diffStage_counterOnePixelStream_payload);
  always @(*) begin
    diffStage_counterOnePixelStream_s2mPipe_ready = resultStage_counterOnePixelStream_ready;
    if(when_Stream_l368_27) begin
      diffStage_counterOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_27 = (! resultStage_counterOnePixelStream_valid);
  assign resultStage_counterOnePixelStream_valid = diffStage_counterOnePixelStream_s2mPipe_rValid;
  assign resultStage_counterOnePixelStream_payload = diffStage_counterOnePixelStream_s2mPipe_rData;
  assign diffStage_mainTwoPixelStream_ready = (! diffStage_mainTwoPixelStream_rValid);
  assign diffStage_mainTwoPixelStream_s2mPipe_valid = (diffStage_mainTwoPixelStream_valid || diffStage_mainTwoPixelStream_rValid);
  assign diffStage_mainTwoPixelStream_s2mPipe_payload = (diffStage_mainTwoPixelStream_rValid ? diffStage_mainTwoPixelStream_rData : diffStage_mainTwoPixelStream_payload);
  always @(*) begin
    diffStage_mainTwoPixelStream_s2mPipe_ready = resultStage_mainTwoPixelStream_ready;
    if(when_Stream_l368_28) begin
      diffStage_mainTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_28 = (! resultStage_mainTwoPixelStream_valid);
  assign resultStage_mainTwoPixelStream_valid = diffStage_mainTwoPixelStream_s2mPipe_rValid;
  assign resultStage_mainTwoPixelStream_payload = diffStage_mainTwoPixelStream_s2mPipe_rData;
  assign diffStage_counterTwoPixelStream_ready = (! diffStage_counterTwoPixelStream_rValid);
  assign diffStage_counterTwoPixelStream_s2mPipe_valid = (diffStage_counterTwoPixelStream_valid || diffStage_counterTwoPixelStream_rValid);
  assign diffStage_counterTwoPixelStream_s2mPipe_payload = (diffStage_counterTwoPixelStream_rValid ? diffStage_counterTwoPixelStream_rData : diffStage_counterTwoPixelStream_payload);
  always @(*) begin
    diffStage_counterTwoPixelStream_s2mPipe_ready = resultStage_counterTwoPixelStream_ready;
    if(when_Stream_l368_29) begin
      diffStage_counterTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_29 = (! resultStage_counterTwoPixelStream_valid);
  assign resultStage_counterTwoPixelStream_valid = diffStage_counterTwoPixelStream_s2mPipe_rValid;
  assign resultStage_counterTwoPixelStream_payload = diffStage_counterTwoPixelStream_s2mPipe_rData;
  assign diffStage_oddRowPixelStream_ready = (! diffStage_oddRowPixelStream_rValid);
  assign diffStage_oddRowPixelStream_s2mPipe_valid = (diffStage_oddRowPixelStream_valid || diffStage_oddRowPixelStream_rValid);
  assign diffStage_oddRowPixelStream_s2mPipe_payload = (diffStage_oddRowPixelStream_rValid ? diffStage_oddRowPixelStream_rData : diffStage_oddRowPixelStream_payload);
  always @(*) begin
    diffStage_oddRowPixelStream_s2mPipe_ready = resultStage_oddRowPixelStream_ready;
    if(when_Stream_l368_30) begin
      diffStage_oddRowPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_30 = (! resultStage_oddRowPixelStream_valid);
  assign resultStage_oddRowPixelStream_valid = diffStage_oddRowPixelStream_s2mPipe_rValid;
  assign resultStage_oddRowPixelStream_payload = diffStage_oddRowPixelStream_s2mPipe_rData;
  assign diffStage_controlPipe_ready = diffStage_controlPipe_fork_io_input_ready;
  assign CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceMode = diffStage_controlPipe_payload_onceMode;
  assign CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceValid = diffStage_controlPipe_payload_onceValid;
  assign CICC1851_when_SuperResolutionPart2_l419 = diffStage_controlPipe_payload_mainDiff;
  assign CICC1851_when_SuperResolutionPart2_l428 = diffStage_controlPipe_payload_counterDiff;
  assign CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceCompValid = diffStage_controlPipe_payload_twiceCompValid;
  assign CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceMode = diffStage_controlPipe_payload_twiceMode;
  always @(*) begin
    CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag = diffStage_controlPipe_payload_inpValidFlag;
    if(CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceValid) begin
      case(CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceMode)
        3'b000 : begin
          if(when_SuperResolutionPart2_l419) begin
            CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag = 1'b0;
          end
        end
        3'b001 : begin
          if(when_SuperResolutionPart2_l420) begin
            CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag = 1'b0;
          end
        end
        3'b010 : begin
          if(when_SuperResolutionPart2_l421) begin
            CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag = 1'b0;
          end
        end
        3'b011 : begin
          if(when_SuperResolutionPart2_l422) begin
            CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag = 1'b0;
          end
        end
        default : begin
        end
      endcase
    end
    if(CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceCompValid) begin
      case(CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceMode)
        3'b000 : begin
          if(when_SuperResolutionPart2_l428) begin
            CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag = 1'b0;
          end
        end
        3'b001 : begin
          if(when_SuperResolutionPart2_l429) begin
            CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag = 1'b0;
          end
        end
        3'b011 : begin
          if(when_SuperResolutionPart2_l430) begin
            CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag = 1'b0;
          end
        end
        3'b101 : begin
          if(when_SuperResolutionPart2_l431) begin
            CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag = 1'b0;
          end
        end
        default : begin
        end
      endcase
    end
  end

  assign when_SuperResolutionPart2_l419 = (inpThreshold <= CICC1851_when_SuperResolutionPart2_l419);
  assign when_SuperResolutionPart2_l420 = (inpThreshold <= CICC1851_when_SuperResolutionPart2_l419);
  assign when_SuperResolutionPart2_l421 = (inpThreshold <= CICC1851_when_SuperResolutionPart2_l419);
  assign when_SuperResolutionPart2_l422 = (inpThreshold <= CICC1851_when_SuperResolutionPart2_l419);
  assign when_SuperResolutionPart2_l428 = ((inpThreshold <= CICC1851_when_SuperResolutionPart2_l419) && (inpThreshold <= CICC1851_when_SuperResolutionPart2_l428));
  assign when_SuperResolutionPart2_l429 = ((inpThreshold <= CICC1851_when_SuperResolutionPart2_l419) && (inpThreshold <= CICC1851_when_SuperResolutionPart2_l428));
  assign when_SuperResolutionPart2_l430 = (inpThreshold <= CICC1851_when_SuperResolutionPart2_l419);
  assign when_SuperResolutionPart2_l431 = (inpThreshold <= CICC1851_when_SuperResolutionPart2_l419);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_valid = diffStage_controlPipe_fork_io_outputs_0_valid;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_payload_frameStart = diffStage_controlPipe_payload_frameStart;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_payload_rowEnd = diffStage_controlPipe_payload_rowEnd;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_payload_passMode = diffStage_controlPipe_payload_passMode;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_payload_passValid = diffStage_controlPipe_payload_passValid;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceMode = CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceMode;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceValid = CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceValid;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_payload_mainCompare = diffStage_controlPipe_payload_mainCompare;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_payload_counterCompare = diffStage_controlPipe_payload_counterCompare;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_payload_mainDiff = CICC1851_when_SuperResolutionPart2_l419;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_payload_counterDiff = CICC1851_when_SuperResolutionPart2_l428;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceCompValid = CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceCompValid;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceMode = CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceMode;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag = CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_payload_oddValid = diffStage_controlPipe_payload_oddValid;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_ready = (! diffStage_controlPipe_fork_io_outputs_0_translated_rValid);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_valid = (diffStage_controlPipe_fork_io_outputs_0_translated_valid || diffStage_controlPipe_fork_io_outputs_0_translated_rValid);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_frameStart = (diffStage_controlPipe_fork_io_outputs_0_translated_rValid ? diffStage_controlPipe_fork_io_outputs_0_translated_rData_frameStart : diffStage_controlPipe_fork_io_outputs_0_translated_payload_frameStart);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_rowEnd = (diffStage_controlPipe_fork_io_outputs_0_translated_rValid ? diffStage_controlPipe_fork_io_outputs_0_translated_rData_rowEnd : diffStage_controlPipe_fork_io_outputs_0_translated_payload_rowEnd);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_passMode = (diffStage_controlPipe_fork_io_outputs_0_translated_rValid ? diffStage_controlPipe_fork_io_outputs_0_translated_rData_passMode : diffStage_controlPipe_fork_io_outputs_0_translated_payload_passMode);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_passValid = (diffStage_controlPipe_fork_io_outputs_0_translated_rValid ? diffStage_controlPipe_fork_io_outputs_0_translated_rData_passValid : diffStage_controlPipe_fork_io_outputs_0_translated_payload_passValid);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_onceMode = (diffStage_controlPipe_fork_io_outputs_0_translated_rValid ? diffStage_controlPipe_fork_io_outputs_0_translated_rData_onceMode : diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceMode);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_onceValid = (diffStage_controlPipe_fork_io_outputs_0_translated_rValid ? diffStage_controlPipe_fork_io_outputs_0_translated_rData_onceValid : diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceValid);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_mainCompare = (diffStage_controlPipe_fork_io_outputs_0_translated_rValid ? diffStage_controlPipe_fork_io_outputs_0_translated_rData_mainCompare : diffStage_controlPipe_fork_io_outputs_0_translated_payload_mainCompare);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_counterCompare = (diffStage_controlPipe_fork_io_outputs_0_translated_rValid ? diffStage_controlPipe_fork_io_outputs_0_translated_rData_counterCompare : diffStage_controlPipe_fork_io_outputs_0_translated_payload_counterCompare);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_mainDiff = (diffStage_controlPipe_fork_io_outputs_0_translated_rValid ? diffStage_controlPipe_fork_io_outputs_0_translated_rData_mainDiff : diffStage_controlPipe_fork_io_outputs_0_translated_payload_mainDiff);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_counterDiff = (diffStage_controlPipe_fork_io_outputs_0_translated_rValid ? diffStage_controlPipe_fork_io_outputs_0_translated_rData_counterDiff : diffStage_controlPipe_fork_io_outputs_0_translated_payload_counterDiff);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_twiceCompValid = (diffStage_controlPipe_fork_io_outputs_0_translated_rValid ? diffStage_controlPipe_fork_io_outputs_0_translated_rData_twiceCompValid : diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceCompValid);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_twiceMode = (diffStage_controlPipe_fork_io_outputs_0_translated_rValid ? diffStage_controlPipe_fork_io_outputs_0_translated_rData_twiceMode : diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceMode);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_inpValidFlag = (diffStage_controlPipe_fork_io_outputs_0_translated_rValid ? diffStage_controlPipe_fork_io_outputs_0_translated_rData_inpValidFlag : diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_oddValid = (diffStage_controlPipe_fork_io_outputs_0_translated_rValid ? diffStage_controlPipe_fork_io_outputs_0_translated_rData_oddValid : diffStage_controlPipe_fork_io_outputs_0_translated_payload_oddValid);
  always @(*) begin
    diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_ready = resultStage_controlPipe_ready;
    if(when_Stream_l368_31) begin
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_31 = (! resultStage_controlPipe_valid);
  assign resultStage_controlPipe_valid = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rValid;
  assign resultStage_controlPipe_payload_frameStart = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_frameStart;
  assign resultStage_controlPipe_payload_rowEnd = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_rowEnd;
  assign resultStage_controlPipe_payload_passMode = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_passMode;
  assign resultStage_controlPipe_payload_passValid = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_passValid;
  assign resultStage_controlPipe_payload_onceMode = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_onceMode;
  assign resultStage_controlPipe_payload_onceValid = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_onceValid;
  assign resultStage_controlPipe_payload_mainCompare = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_mainCompare;
  assign resultStage_controlPipe_payload_counterCompare = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_counterCompare;
  assign resultStage_controlPipe_payload_mainDiff = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_mainDiff;
  assign resultStage_controlPipe_payload_counterDiff = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_counterDiff;
  assign resultStage_controlPipe_payload_twiceCompValid = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_twiceCompValid;
  assign resultStage_controlPipe_payload_twiceMode = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_twiceMode;
  assign resultStage_controlPipe_payload_inpValidFlag = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_inpValidFlag;
  assign resultStage_controlPipe_payload_oddValid = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_oddValid;
  assign resultStage_pixelStream_valid = diffStage_controlPipe_fork_io_outputs_1_valid;
  always @(*) begin
    resultStage_pixelStream_payload = 8'h0;
    if(diffStage_controlPipe_fork_io_outputs_1_payload_passValid) begin
      if(diffStage_controlPipe_fork_io_outputs_1_payload_passMode) begin
        resultStage_pixelStream_payload = diffStage_mainTwoPixelStream_payload;
      end else begin
        resultStage_pixelStream_payload = diffStage_mainOnePixelStream_payload;
      end
    end
    if(diffStage_controlPipe_fork_io_outputs_1_payload_oddValid) begin
      resultStage_pixelStream_payload = diffStage_oddRowPixelStream_payload;
    end
    if(diffStage_controlPipe_fork_io_outputs_1_payload_onceValid) begin
      case(diffStage_controlPipe_fork_io_outputs_1_payload_onceMode)
        3'b000 : begin
          if(when_SuperResolutionPart2_l451) begin
            resultStage_pixelStream_payload = 8'h0;
          end else begin
            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload[7:0];
          end
        end
        3'b001 : begin
          if(when_SuperResolutionPart2_l455) begin
            resultStage_pixelStream_payload = 8'h0;
          end else begin
            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_2[7:0];
          end
        end
        3'b010 : begin
          if(when_SuperResolutionPart2_l459) begin
            resultStage_pixelStream_payload = 8'h0;
          end else begin
            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_4[7:0];
          end
        end
        3'b011 : begin
          if(when_SuperResolutionPart2_l463) begin
            resultStage_pixelStream_payload = 8'h0;
          end else begin
            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_6[7:0];
          end
        end
        3'b100 : begin
          resultStage_pixelStream_payload = diffStage_mainOnePixelStream_payload;
        end
        3'b101 : begin
          resultStage_pixelStream_payload = diffStage_mainTwoPixelStream_payload;
        end
        default : begin
        end
      endcase
    end
    if(diffStage_controlPipe_fork_io_outputs_1_payload_twiceCompValid) begin
      case(diffStage_controlPipe_fork_io_outputs_1_payload_twiceMode)
        3'b000 : begin
          if(when_SuperResolutionPart2_l474) begin
            resultStage_pixelStream_payload = 8'h0;
          end else begin
            if(when_SuperResolutionPart2_l477) begin
              resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_8[7:0];
            end else begin
              resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_10[7:0];
            end
          end
        end
        3'b001 : begin
          if(when_SuperResolutionPart2_l482) begin
            resultStage_pixelStream_payload = 8'h0;
          end else begin
            if(when_SuperResolutionPart2_l485) begin
              resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_12[7:0];
            end else begin
              resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_14[7:0];
            end
          end
        end
        3'b010 : begin
          resultStage_pixelStream_payload = diffStage_mainTwoPixelStream_payload;
        end
        3'b011 : begin
          if(when_SuperResolutionPart2_l491) begin
            resultStage_pixelStream_payload = 8'h0;
          end else begin
            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_16[7:0];
          end
        end
        3'b100 : begin
          resultStage_pixelStream_payload = diffStage_mainOnePixelStream_payload;
        end
        3'b101 : begin
          if(when_SuperResolutionPart2_l496) begin
            resultStage_pixelStream_payload = 8'h0;
          end else begin
            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_18[7:0];
          end
        end
        default : begin
        end
      endcase
    end
  end

  assign when_SuperResolutionPart2_l451 = (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart2_l455 = (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart2_l459 = (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart2_l463 = (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart2_l474 = ((inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff) && (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff));
  assign when_SuperResolutionPart2_l477 = (diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart2_l482 = ((inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff) && (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff));
  assign when_SuperResolutionPart2_l485 = (diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart2_l491 = (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart2_l496 = (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign resultStage_pixelStream_ready = (! resultStage_pixelStream_rValid);
  assign resultStage_pixelStream_s2mPipe_valid = (resultStage_pixelStream_valid || resultStage_pixelStream_rValid);
  assign resultStage_pixelStream_s2mPipe_payload = (resultStage_pixelStream_rValid ? resultStage_pixelStream_rData : resultStage_pixelStream_payload);
  always @(*) begin
    resultStage_pixelStream_s2mPipe_ready = resultStage_resultStream_ready;
    if(when_Stream_l368_32) begin
      resultStage_pixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_32 = (! resultStage_resultStream_valid);
  assign resultStage_resultStream_valid = resultStage_pixelStream_s2mPipe_rValid;
  assign resultStage_resultStream_payload = resultStage_pixelStream_s2mPipe_rData;
  assign CICC1851_resultStage_mainOnePixelStream_ready_2 = (CICC1851_resultStage_mainOnePixelStream_ready && CICC1851_resultStage_mainOnePixelStream_ready_1);
  assign CICC1851_resultStage_mainOnePixelStream_ready = ((((((resultStage_resultStream_valid && resultStage_mainOnePixelStream_valid) && resultStage_counterOnePixelStream_valid) && resultStage_mainTwoPixelStream_valid) && resultStage_counterTwoPixelStream_valid) && resultStage_controlPipe_valid) && resultStage_oddRowPixelStream_valid);
  assign resultStage_resultStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_mainOnePixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_counterOnePixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_mainTwoPixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_counterTwoPixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_controlPipe_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_oddRowPixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign when_Stream_l438 = ((((! resultStage_controlPipe_payload_passValid) && (! resultStage_controlPipe_payload_onceValid)) && (! resultStage_controlPipe_payload_twiceCompValid)) && (! resultStage_controlPipe_payload_oddValid));
  always @(*) begin
    resultsJoin_valid = CICC1851_resultStage_mainOnePixelStream_ready;
    if(when_Stream_l438) begin
      resultsJoin_valid = 1'b0;
    end
  end

  always @(*) begin
    CICC1851_resultStage_mainOnePixelStream_ready_1 = resultsJoin_ready;
    if(when_Stream_l438) begin
      CICC1851_resultStage_mainOnePixelStream_ready_1 = 1'b1;
    end
  end

  assign pixelsStream_valid = resultsJoin_valid;
  assign resultsJoin_ready = pixelsStream_ready;
  assign pixelsStream_payload_pixel = resultStage_resultStream_payload;
  assign pixelsStream_payload_frameStart = resultStage_controlPipe_payload_frameStart;
  assign pixelsStream_payload_rowEnd = resultStage_controlPipe_payload_rowEnd;
  assign pixelsStream_payload_inpValid = resultStage_controlPipe_payload_inpValidFlag;
  assign pixelsStream_ready = (! pixelsStream_rValid);
  assign pixelsStream_s2mPipe_valid = (pixelsStream_valid || pixelsStream_rValid);
  assign pixelsStream_s2mPipe_payload_pixel = (pixelsStream_rValid ? pixelsStream_rData_pixel : pixelsStream_payload_pixel);
  assign pixelsStream_s2mPipe_payload_frameStart = (pixelsStream_rValid ? pixelsStream_rData_frameStart : pixelsStream_payload_frameStart);
  assign pixelsStream_s2mPipe_payload_rowEnd = (pixelsStream_rValid ? pixelsStream_rData_rowEnd : pixelsStream_payload_rowEnd);
  assign pixelsStream_s2mPipe_payload_inpValid = (pixelsStream_rValid ? pixelsStream_rData_inpValid : pixelsStream_payload_inpValid);
  always @(*) begin
    pixelsStream_s2mPipe_ready = pixelsStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_33) begin
      pixelsStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_33 = (! pixelsStream_s2mPipe_m2sPipe_valid);
  assign pixelsStream_s2mPipe_m2sPipe_valid = pixelsStream_s2mPipe_rValid;
  assign pixelsStream_s2mPipe_m2sPipe_payload_pixel = pixelsStream_s2mPipe_rData_pixel;
  assign pixelsStream_s2mPipe_m2sPipe_payload_frameStart = pixelsStream_s2mPipe_rData_frameStart;
  assign pixelsStream_s2mPipe_m2sPipe_payload_rowEnd = pixelsStream_s2mPipe_rData_rowEnd;
  assign pixelsStream_s2mPipe_m2sPipe_payload_inpValid = pixelsStream_s2mPipe_rData_inpValid;
  assign pixelsStream_s2mPipe_m2sPipe_ready = pixelsOut_ready;
  assign controlStateMachine_wantExit = 1'b0;
  always @(*) begin
    controlStateMachine_wantStart = 1'b0;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_4_HOLD : begin
      end
      controlStateMachine_enumDef_4_PASS : begin
      end
      controlStateMachine_enumDef_4_ONCE : begin
      end
      controlStateMachine_enumDef_4_TWICE : begin
      end
      default : begin
        controlStateMachine_wantStart = 1'b1;
      end
    endcase
  end

  assign controlStateMachine_wantKill = 1'b0;
  assign when_SuperResolutionPart2_l761 = (((currentState == 3'b010) || (currentState == 3'b011)) || (currentState == 3'b100));
  assign controlStream_fire_4 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart2_l763 = (controlStream_fire_4 && (CICC1851_when_SuperResolutionPart2_l763 == CICC1851_when_SuperResolutionPart2_l763_1));
  assign controlStream_fire_5 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart2_l764 = ((outReachRowEnd && (CICC1851_when_SuperResolutionPart2_l764 == CICC1851_when_SuperResolutionPart2_l764_1)) && controlStream_fire_5);
  assign controlStream_fire_6 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart2_l766 = (controlStream_fire_6 && outReachRowEnd);
  assign controlStream_fire_7 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart2_l783 = (CICC1851_when_SuperResolutionPart2_l783 == 12'h0);
  assign when_SuperResolutionPart2_l785 = (CICC1851_when_SuperResolutionPart2_l785 == 12'h001);
  assign when_SuperResolutionPart2_l787 = (CICC1851_when_SuperResolutionPart2_l787 == 12'h002);
  assign when_SuperResolutionPart2_l789 = (CICC1851_when_SuperResolutionPart2_l789 == 12'h003);
  assign when_SuperResolutionPart2_l793 = (CICC1851_when_SuperResolutionPart2_l793 == 12'h0);
  assign when_SuperResolutionPart2_l796 = (CICC1851_when_SuperResolutionPart2_l796 == 12'h001);
  assign when_SuperResolutionPart2_l799 = (CICC1851_when_SuperResolutionPart2_l799 == 12'h002);
  assign when_SuperResolutionPart2_l802 = (CICC1851_when_SuperResolutionPart2_l802 == 12'h003);
  always @(*) begin
    controlStateMachine_stateNext = controlStateMachine_stateReg;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_4_HOLD : begin
        if(zeroInFourOutRow) begin
          if(passPixels_fire_13) begin
            if(threeInFourOutPixelAddr) begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_4_ONCE;
            end else begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_4_PASS;
            end
          end
        end else begin
          if(twoInFourOutRow) begin
            if(passPixels_fire_14) begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_4_PASS;
            end
          end else begin
            if(threeInFourOutRow) begin
              if(passPixels_fire_15) begin
                if(threeInFourOutPixelAddr) begin
                  if(willHoldToTwice) begin
                    controlStateMachine_stateNext = controlStateMachine_enumDef_4_TWICE;
                  end
                end else begin
                  controlStateMachine_stateNext = controlStateMachine_enumDef_4_ONCE;
                end
              end
            end
          end
        end
      end
      controlStateMachine_enumDef_4_PASS : begin
        if(controlStream_fire_8) begin
          if(oneInFourOutPixelAddr) begin
            if(oneInFourOutRow) begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_4_PASS;
            end else begin
              if(twoInFourOutRow) begin
                if(when_SuperResolutionPart2_l573) begin
                  controlStateMachine_stateNext = controlStateMachine_enumDef_4_HOLD;
                end else begin
                  controlStateMachine_stateNext = controlStateMachine_enumDef_4_PASS;
                end
              end else begin
                if(when_SuperResolutionPart2_l578) begin
                  controlStateMachine_stateNext = controlStateMachine_enumDef_4_HOLD;
                end else begin
                  controlStateMachine_stateNext = controlStateMachine_enumDef_4_PASS;
                end
              end
            end
          end else begin
            if(twoInFourOutPixelAddr) begin
              if(oneInFourOutRow) begin
                controlStateMachine_stateNext = controlStateMachine_enumDef_4_ONCE;
              end else begin
                if(twoInFourOutRow) begin
                  controlStateMachine_stateNext = controlStateMachine_enumDef_4_ONCE;
                end else begin
                  if(when_SuperResolutionPart2_l590) begin
                    controlStateMachine_stateNext = controlStateMachine_enumDef_4_HOLD;
                  end else begin
                    controlStateMachine_stateNext = controlStateMachine_enumDef_4_ONCE;
                  end
                end
              end
            end else begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_4_PASS;
            end
          end
        end
      end
      controlStateMachine_enumDef_4_ONCE : begin
        if(controlStream_fire_10) begin
          if(zeroInFourOutRow) begin
            controlStateMachine_stateNext = controlStateMachine_enumDef_4_PASS;
          end else begin
            if(oneInFourOutRow) begin
              if(when_SuperResolutionPart2_l642) begin
                controlStateMachine_stateNext = controlStateMachine_enumDef_4_HOLD;
              end else begin
                controlStateMachine_stateNext = controlStateMachine_enumDef_4_PASS;
              end
            end else begin
              if(twoInFourOutRow) begin
                if(outReachRowEnd) begin
                  if(when_SuperResolutionPart2_l647) begin
                    controlStateMachine_stateNext = controlStateMachine_enumDef_4_HOLD;
                  end else begin
                    controlStateMachine_stateNext = controlStateMachine_enumDef_4_ONCE;
                  end
                end else begin
                  controlStateMachine_stateNext = controlStateMachine_enumDef_4_PASS;
                end
              end else begin
                if(twoInFourOutPixelAddr) begin
                  if(when_SuperResolutionPart2_l653) begin
                    controlStateMachine_stateNext = controlStateMachine_enumDef_4_HOLD;
                  end else begin
                    controlStateMachine_stateNext = controlStateMachine_enumDef_4_TWICE;
                  end
                end else begin
                  controlStateMachine_stateNext = controlStateMachine_enumDef_4_ONCE;
                end
              end
            end
          end
        end
      end
      controlStateMachine_enumDef_4_TWICE : begin
        if(controlStream_fire_11) begin
          if(outReachRowEnd) begin
            if(outReachFinalRow) begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_4_HOLD;
            end else begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_4_PASS;
            end
          end else begin
            controlStateMachine_stateNext = controlStateMachine_enumDef_4_ONCE;
          end
        end
      end
      default : begin
      end
    endcase
    if(controlStateMachine_wantStart) begin
      controlStateMachine_stateNext = controlStateMachine_enumDef_4_HOLD;
    end
    if(controlStateMachine_wantKill) begin
      controlStateMachine_stateNext = controlStateMachine_enumDef_4_BOOT;
    end
  end

  assign passPixels_fire_13 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_14 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_15 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_16 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart2_l560 = (CICC1851_when_SuperResolutionPart2_l560 == CICC1851_when_SuperResolutionPart2_l560_1);
  assign controlStream_fire_8 = (controlStream_valid && controlStream_ready);
  assign passPixels_fire_17 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart2_l573 = ((((oddBufferRow && (! holdBuffer)) && willPassToHoldCaseOne) && (! passPixels_fire_17)) && (! bufferReuse));
  assign passPixels_fire_18 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart2_l578 = (((((! oddBufferRow) && (! holdBuffer)) && willPassToHoldCaseOne) && (! passPixels_fire_18)) && (! bufferReuse));
  assign when_SuperResolutionPart2_l585 = ((oddBufferRow && (! holdBuffer)) && (! bufferReachRowEnd));
  assign when_SuperResolutionPart2_l588 = (((! oddBufferRow) && (! bufferReuse)) && (! bufferReachRowEnd));
  assign passPixels_fire_19 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart2_l590 = (((((! oddBufferRow) && (! holdBuffer)) && (! bufferReuse)) && (willPassToHoldCaseTwo || holdWillPassToHoldCaseTwo)) && (! passPixels_fire_19));
  assign when_SuperResolutionPart2_l602 = (poping && (CICC1851_when_SuperResolutionPart2_l602 == CICC1851_when_SuperResolutionPart2_l602_1));
  assign when_SuperResolutionPart2_l603 = (pushAndPoping && (CICC1851_when_SuperResolutionPart2_l603 == CICC1851_when_SuperResolutionPart2_l603_1));
  assign when_SuperResolutionPart2_l605 = (poping && (CICC1851_when_SuperResolutionPart2_l605 == CICC1851_when_SuperResolutionPart2_l605_1));
  assign when_SuperResolutionPart2_l606 = (pushAndPoping && (CICC1851_when_SuperResolutionPart2_l606 == CICC1851_when_SuperResolutionPart2_l606_1));
  assign when_SuperResolutionPart2_l609 = (CICC1851_when_SuperResolutionPart2_l609 == 12'h0);
  assign controlStream_fire_9 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart2_l630 = (frameStart && controlStream_fire_9);
  assign controlStream_fire_10 = (controlStream_valid && controlStream_ready);
  assign passPixels_fire_20 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart2_l642 = (((outReachRowEnd && willOnceToHoldCaseOne) && (bufferWAddr_value == 11'h0)) && (! passPixels_fire_20));
  assign passPixels_fire_21 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart2_l647 = (((bufferWAddr_value == 11'h0) && (! passPixels_fire_21)) && willOnceToHoldCaseTwo);
  assign passPixels_fire_22 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart2_l653 = ((((! oddBufferRow) && willOnceToHoldCaseThree) && (! passPixels_fire_22)) && (! bufferReuse));
  assign passPixels_fire_23 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart2_l662 = (passPixels_fire_23 && bufferReachRowEnd);
  assign when_SuperResolutionPart2_l667 = (poping && (CICC1851_when_SuperResolutionPart2_l667 == CICC1851_when_SuperResolutionPart2_l667_2));
  assign when_SuperResolutionPart2_l668 = (pushAndPoping && (CICC1851_when_SuperResolutionPart2_l668 == CICC1851_when_SuperResolutionPart2_l668_1));
  assign controlStream_fire_11 = (controlStream_valid && controlStream_ready);
  assign currentState = controlStateMachine_stateReg;
  always @(posedge clk or negedge resetn) begin
    if(!resetn) begin
      inpTwoDone <= 1'b0;
      readDone <= 1'b0;
      startRead <= 1'b0;
      slaveStart <= 1'b0;
      frameStart <= 1'b0;
      inpThreshold <= 8'h80;
      bmpWidth <= 10'h3c0;
      bmpHeight <= 10'h21c;
      holdBuffer <= 1'b0;
      writeDone <= 1'b0;
      bufferRowCount_value <= 11'h0;
      bufferReuse <= 1'b0;
      bufferEnable <= 1'b0;
      bufferSwitch <= 2'b00;
      nextRowBuffer <= 1'b1;
      bufferWAddr_value <= 11'h0;
      outPixelAddr_value <= 12'h0;
      outRowCount_value <= 12'h0;
      alreadySendRow_value <= 12'h0;
      alreadySendCountInRow_value <= 12'h0;
      alreadyReachRowEnd <= 1'b0;
      alreadyReachFinalRow <= 1'b0;
      outReachRowEnd <= 1'b0;
      outReachFinalRow <= 1'b0;
      bufferReachRowEnd <= 1'b0;
      bufferReachFinalRow <= 1'b0;
      oddBufferRow <= 1'b0;
      zeroInFourOutPixelAddr <= 1'b1;
      oneInFourOutPixelAddr <= 1'b0;
      twoInFourOutPixelAddr <= 1'b0;
      threeInFourOutPixelAddr <= 1'b0;
      zeroInFourOutRow <= 1'b1;
      oneInFourOutRow <= 1'b0;
      twoInFourOutRow <= 1'b0;
      threeInFourOutRow <= 1'b0;
      willHoldToTwice <= 1'b0;
      willPassToHoldCaseOne <= 1'b0;
      willPassToHoldCaseTwo <= 1'b0;
      holdWillPassToHoldCaseTwo <= 1'b0;
      willOnceToHoldCaseOne <= 1'b0;
      willOnceToHoldCaseTwo <= 1'b0;
      willOnceToHoldCaseThree <= 1'b0;
      pixelsIn_rValid <= 1'b0;
      pixelsIn_s2mPipe_rValid <= 1'b0;
      mainAddrOneStream_rValid <= 1'b0;
      mainAddrOneStream_s2mPipe_rValid <= 1'b0;
      CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_mainOnePixelStream_valid <= 1'b0;
      counterAddrOneStream_rValid <= 1'b0;
      counterAddrOneStream_s2mPipe_rValid <= 1'b0;
      CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_counterOnePixelStream_valid <= 1'b0;
      mainAddrTwoStream_rValid <= 1'b0;
      mainAddrTwoStream_s2mPipe_rValid <= 1'b0;
      CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_mainTwoPixelStream_valid <= 1'b0;
      counterAddrTwoStream_rValid <= 1'b0;
      counterAddrTwoStream_s2mPipe_rValid <= 1'b0;
      CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_counterTwoPixelStream_valid <= 1'b0;
      oddAddrStream_rValid <= 1'b0;
      oddAddrStream_s2mPipe_rValid <= 1'b0;
      CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_oddRowPixelStream_valid <= 1'b0;
      controlStream_rValid <= 1'b0;
      controlStream_s2mPipe_rValid <= 1'b0;
      controlStream_s2mPipe_m2sPipe_rValid <= 1'b0;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rValid <= 1'b0;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rValid <= 1'b0;
      readStage_mainOnePixelStream_rValid <= 1'b0;
      readStage_mainOnePixelStream_s2mPipe_rValid <= 1'b0;
      readStage_counterOnePixelStream_rValid <= 1'b0;
      readStage_counterOnePixelStream_s2mPipe_rValid <= 1'b0;
      readStage_mainTwoPixelStream_rValid <= 1'b0;
      readStage_mainTwoPixelStream_s2mPipe_rValid <= 1'b0;
      readStage_counterTwoPixelStream_rValid <= 1'b0;
      readStage_counterTwoPixelStream_s2mPipe_rValid <= 1'b0;
      readStage_oddRowPixelStream_rValid <= 1'b0;
      readStage_oddRowPixelStream_s2mPipe_rValid <= 1'b0;
      readStage_controlPipe_translated_rValid <= 1'b0;
      readStage_controlPipe_translated_s2mPipe_rValid <= 1'b0;
      compareStage_mainOnePixelStream_rValid <= 1'b0;
      compareStage_mainOnePixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_counterOnePixelStream_rValid <= 1'b0;
      compareStage_counterOnePixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_mainTwoPixelStream_rValid <= 1'b0;
      compareStage_mainTwoPixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_counterTwoPixelStream_rValid <= 1'b0;
      compareStage_counterTwoPixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_oddRowPixelStream_rValid <= 1'b0;
      compareStage_oddRowPixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_controlPipe_translated_rValid <= 1'b0;
      compareStage_controlPipe_translated_s2mPipe_rValid <= 1'b0;
      diffStage_mainOnePixelStream_rValid <= 1'b0;
      diffStage_mainOnePixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_counterOnePixelStream_rValid <= 1'b0;
      diffStage_counterOnePixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_mainTwoPixelStream_rValid <= 1'b0;
      diffStage_mainTwoPixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_counterTwoPixelStream_rValid <= 1'b0;
      diffStage_counterTwoPixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_oddRowPixelStream_rValid <= 1'b0;
      diffStage_oddRowPixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_controlPipe_fork_io_outputs_0_translated_rValid <= 1'b0;
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rValid <= 1'b0;
      resultStage_pixelStream_rValid <= 1'b0;
      resultStage_pixelStream_s2mPipe_rValid <= 1'b0;
      pixelsStream_rValid <= 1'b0;
      pixelsStream_s2mPipe_rValid <= 1'b0;
      controlStateMachine_stateReg <= controlStateMachine_enumDef_4_BOOT;
    end else begin
      if(when_SuperResolutionPart2_l40) begin
        inpTwoDone <= 1'b0;
      end
      if(when_SuperResolutionPart2_l43) begin
        readDone <= 1'b0;
      end
      if(when_SuperResolutionPart2_l46) begin
        startRead <= 1'b1;
      end
      if(when_SuperResolutionPart2_l46_1) begin
        startRead <= 1'b0;
      end
      if(when_SuperResolutionPart2_l49) begin
        slaveStart <= 1'b1;
      end
      if(when_SuperResolutionPart2_l49_1) begin
        slaveStart <= 1'b0;
      end
      inpThreshold <= thresholdIn;
      bmpWidth <= widthIn;
      bmpHeight <= heightIn;
      if(when_SuperResolutionPart2_l64) begin
        holdBuffer <= 1'b0;
      end
      if(when_SuperResolutionPart2_l67) begin
        writeDone <= 1'b0;
      end
      bufferRowCount_value <= bufferRowCount_valueNext;
      if(inpTwoDone) begin
        bufferReuse <= 1'b0;
      end
      if(when_SuperResolutionPart2_l76) begin
        bufferEnable <= 1'b1;
      end
      if(when_SuperResolutionPart2_l76_1) begin
        bufferEnable <= 1'b0;
      end
      if(when_SuperResolutionPart2_l82) begin
        nextRowBuffer <= 1'b1;
      end
      bufferWAddr_value <= bufferWAddr_valueNext;
      outPixelAddr_value <= outPixelAddr_valueNext;
      outRowCount_value <= outRowCount_valueNext;
      alreadySendRow_value <= alreadySendRow_valueNext;
      alreadySendCountInRow_value <= alreadySendCountInRow_valueNext;
      if(when_SuperResolutionPart2_l106) begin
        oddBufferRow <= 1'b0;
      end
      if(when_SuperResolutionPart2_l108) begin
        zeroInFourOutPixelAddr <= 1'b1;
      end
      if(when_SuperResolutionPart2_l109) begin
        oneInFourOutPixelAddr <= 1'b0;
      end
      if(when_SuperResolutionPart2_l110) begin
        twoInFourOutPixelAddr <= 1'b0;
      end
      if(when_SuperResolutionPart2_l111) begin
        threeInFourOutPixelAddr <= 1'b0;
      end
      if(when_SuperResolutionPart2_l113) begin
        zeroInFourOutRow <= 1'b1;
      end
      if(when_SuperResolutionPart2_l114) begin
        oneInFourOutRow <= 1'b0;
      end
      if(when_SuperResolutionPart2_l115) begin
        twoInFourOutRow <= 1'b0;
      end
      if(when_SuperResolutionPart2_l116) begin
        threeInFourOutRow <= 1'b0;
      end
      if(when_SuperResolutionPart2_l120) begin
        willHoldToTwice <= 1'b0;
      end
      if(when_SuperResolutionPart2_l121) begin
        willPassToHoldCaseOne <= 1'b0;
      end
      if(when_SuperResolutionPart2_l122) begin
        willPassToHoldCaseTwo <= 1'b0;
      end
      if(when_SuperResolutionPart2_l123) begin
        holdWillPassToHoldCaseTwo <= 1'b0;
      end
      if(when_SuperResolutionPart2_l124) begin
        willOnceToHoldCaseOne <= 1'b0;
      end
      if(when_SuperResolutionPart2_l125) begin
        willOnceToHoldCaseTwo <= 1'b0;
      end
      if(when_SuperResolutionPart2_l126) begin
        willOnceToHoldCaseThree <= 1'b0;
      end
      if(when_SuperResolutionPart2_l134) begin
        bufferSwitch <= 2'b00;
      end
      if(pixelsIn_valid) begin
        pixelsIn_rValid <= 1'b1;
      end
      if(pixelsIn_s2mPipe_ready) begin
        pixelsIn_rValid <= 1'b0;
      end
      if(pixelsIn_s2mPipe_ready) begin
        pixelsIn_s2mPipe_rValid <= pixelsIn_s2mPipe_valid;
      end
      if(when_SuperResolutionPart2_l181) begin
        bufferReachRowEnd <= 1'b1;
      end
      if(when_SuperResolutionPart2_l182) begin
        bufferReachFinalRow <= 1'b1;
      end
      if(when_SuperResolutionPart2_l185) begin
        if(bufferReachFinalRow) begin
          bufferReachRowEnd <= 1'b0;
          bufferReachFinalRow <= 1'b0;
          bufferReuse <= 1'b1;
        end else begin
          bufferReachRowEnd <= 1'b0;
        end
        if(when_SuperResolutionPart2_l195) begin
          oddBufferRow <= 1'b1;
        end else begin
          oddBufferRow <= 1'b0;
        end
      end
      if(when_SuperResolutionPart2_l200) begin
        if(when_SuperResolutionPart2_l201) begin
          bufferSwitch <= 2'b01;
        end else begin
          if(nextRowBuffer) begin
            bufferSwitch <= (bufferSwitch + 2'b01);
          end else begin
            bufferSwitch <= (bufferSwitch - 2'b01);
          end
        end
      end
      if(when_SuperResolutionPart2_l207) begin
        if(when_SuperResolutionPart2_l208) begin
          holdBuffer <= 1'b1;
          bufferEnable <= 1'b0;
        end
        if(when_SuperResolutionPart2_l212) begin
          writeDone <= 1'b1;
          bufferEnable <= 1'b0;
        end
      end
      if(when_SuperResolutionPart2_l218) begin
        holdBuffer <= 1'b0;
        if(when_SuperResolutionPart2_l220) begin
          nextRowBuffer <= (! nextRowBuffer);
        end
      end
      if(when_SuperResolutionPart2_l224) begin
        frameStart <= 1'b1;
      end
      if(when_SuperResolutionPart2_l234) begin
        alreadyReachRowEnd <= 1'b1;
      end
      if(when_SuperResolutionPart2_l235) begin
        alreadyReachFinalRow <= 1'b1;
      end
      if(pixelsOut_fire_2) begin
        if(alreadyReachRowEnd) begin
          alreadyReachRowEnd <= 1'b0;
          if(alreadyReachFinalRow) begin
            alreadyReachFinalRow <= 1'b0;
          end
        end
      end
      if(when_SuperResolutionPart2_l246) begin
        inpTwoDone <= 1'b1;
      end
      if(mainAddrOneStream_valid) begin
        mainAddrOneStream_rValid <= 1'b1;
      end
      if(mainAddrOneStream_s2mPipe_ready) begin
        mainAddrOneStream_rValid <= 1'b0;
      end
      if(mainAddrOneStream_s2mPipe_ready) begin
        mainAddrOneStream_s2mPipe_rValid <= mainAddrOneStream_s2mPipe_valid;
      end
      if(CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(mainAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_2 <= mainAddrOneStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_1) begin
        CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_1) begin
        CICC1851_readStage_mainOnePixelStream_valid <= (CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready || CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_3);
      end
      if(counterAddrOneStream_valid) begin
        counterAddrOneStream_rValid <= 1'b1;
      end
      if(counterAddrOneStream_s2mPipe_ready) begin
        counterAddrOneStream_rValid <= 1'b0;
      end
      if(counterAddrOneStream_s2mPipe_ready) begin
        counterAddrOneStream_s2mPipe_rValid <= counterAddrOneStream_s2mPipe_valid;
      end
      if(CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(counterAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_2 <= counterAddrOneStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_2) begin
        CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_2) begin
        CICC1851_readStage_counterOnePixelStream_valid <= (CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready || CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_3);
      end
      if(mainAddrTwoStream_valid) begin
        mainAddrTwoStream_rValid <= 1'b1;
      end
      if(mainAddrTwoStream_s2mPipe_ready) begin
        mainAddrTwoStream_rValid <= 1'b0;
      end
      if(mainAddrTwoStream_s2mPipe_ready) begin
        mainAddrTwoStream_s2mPipe_rValid <= mainAddrTwoStream_s2mPipe_valid;
      end
      if(CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(mainAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= mainAddrTwoStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_3) begin
        CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_3) begin
        CICC1851_readStage_mainTwoPixelStream_valid <= (CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready || CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_3);
      end
      if(counterAddrTwoStream_valid) begin
        counterAddrTwoStream_rValid <= 1'b1;
      end
      if(counterAddrTwoStream_s2mPipe_ready) begin
        counterAddrTwoStream_rValid <= 1'b0;
      end
      if(counterAddrTwoStream_s2mPipe_ready) begin
        counterAddrTwoStream_s2mPipe_rValid <= counterAddrTwoStream_s2mPipe_valid;
      end
      if(CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(counterAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= counterAddrTwoStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_4) begin
        CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_4) begin
        CICC1851_readStage_counterTwoPixelStream_valid <= (CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready || CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_3);
      end
      if(oddAddrStream_valid) begin
        oddAddrStream_rValid <= 1'b1;
      end
      if(oddAddrStream_s2mPipe_ready) begin
        oddAddrStream_rValid <= 1'b0;
      end
      if(oddAddrStream_s2mPipe_ready) begin
        oddAddrStream_s2mPipe_rValid <= oddAddrStream_s2mPipe_valid;
      end
      if(CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(oddAddrStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_2 <= oddAddrStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_5) begin
        CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_5) begin
        CICC1851_readStage_oddRowPixelStream_valid <= (CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready || CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_3);
      end
      if(controlStream_valid) begin
        controlStream_rValid <= 1'b1;
      end
      if(controlStream_s2mPipe_ready) begin
        controlStream_rValid <= 1'b0;
      end
      if(controlStream_s2mPipe_ready) begin
        controlStream_s2mPipe_rValid <= controlStream_s2mPipe_valid;
      end
      if(controlStream_s2mPipe_m2sPipe_ready) begin
        controlStream_s2mPipe_m2sPipe_rValid <= controlStream_s2mPipe_m2sPipe_valid;
      end
      if(controlStream_s2mPipe_m2sPipe_m2sPipe_valid) begin
        controlStream_s2mPipe_m2sPipe_m2sPipe_rValid <= 1'b1;
      end
      if(controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready) begin
        controlStream_s2mPipe_m2sPipe_m2sPipe_rValid <= 1'b0;
      end
      if(controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready) begin
        controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_valid;
      end
      if(readStage_mainOnePixelStream_valid) begin
        readStage_mainOnePixelStream_rValid <= 1'b1;
      end
      if(readStage_mainOnePixelStream_s2mPipe_ready) begin
        readStage_mainOnePixelStream_rValid <= 1'b0;
      end
      if(readStage_mainOnePixelStream_s2mPipe_ready) begin
        readStage_mainOnePixelStream_s2mPipe_rValid <= readStage_mainOnePixelStream_s2mPipe_valid;
      end
      if(readStage_counterOnePixelStream_valid) begin
        readStage_counterOnePixelStream_rValid <= 1'b1;
      end
      if(readStage_counterOnePixelStream_s2mPipe_ready) begin
        readStage_counterOnePixelStream_rValid <= 1'b0;
      end
      if(readStage_counterOnePixelStream_s2mPipe_ready) begin
        readStage_counterOnePixelStream_s2mPipe_rValid <= readStage_counterOnePixelStream_s2mPipe_valid;
      end
      if(readStage_mainTwoPixelStream_valid) begin
        readStage_mainTwoPixelStream_rValid <= 1'b1;
      end
      if(readStage_mainTwoPixelStream_s2mPipe_ready) begin
        readStage_mainTwoPixelStream_rValid <= 1'b0;
      end
      if(readStage_mainTwoPixelStream_s2mPipe_ready) begin
        readStage_mainTwoPixelStream_s2mPipe_rValid <= readStage_mainTwoPixelStream_s2mPipe_valid;
      end
      if(readStage_counterTwoPixelStream_valid) begin
        readStage_counterTwoPixelStream_rValid <= 1'b1;
      end
      if(readStage_counterTwoPixelStream_s2mPipe_ready) begin
        readStage_counterTwoPixelStream_rValid <= 1'b0;
      end
      if(readStage_counterTwoPixelStream_s2mPipe_ready) begin
        readStage_counterTwoPixelStream_s2mPipe_rValid <= readStage_counterTwoPixelStream_s2mPipe_valid;
      end
      if(readStage_oddRowPixelStream_valid) begin
        readStage_oddRowPixelStream_rValid <= 1'b1;
      end
      if(readStage_oddRowPixelStream_s2mPipe_ready) begin
        readStage_oddRowPixelStream_rValid <= 1'b0;
      end
      if(readStage_oddRowPixelStream_s2mPipe_ready) begin
        readStage_oddRowPixelStream_s2mPipe_rValid <= readStage_oddRowPixelStream_s2mPipe_valid;
      end
      if(readStage_controlPipe_translated_valid) begin
        readStage_controlPipe_translated_rValid <= 1'b1;
      end
      if(readStage_controlPipe_translated_s2mPipe_ready) begin
        readStage_controlPipe_translated_rValid <= 1'b0;
      end
      if(readStage_controlPipe_translated_s2mPipe_ready) begin
        readStage_controlPipe_translated_s2mPipe_rValid <= readStage_controlPipe_translated_s2mPipe_valid;
      end
      if(compareStage_mainOnePixelStream_valid) begin
        compareStage_mainOnePixelStream_rValid <= 1'b1;
      end
      if(compareStage_mainOnePixelStream_s2mPipe_ready) begin
        compareStage_mainOnePixelStream_rValid <= 1'b0;
      end
      if(compareStage_mainOnePixelStream_s2mPipe_ready) begin
        compareStage_mainOnePixelStream_s2mPipe_rValid <= compareStage_mainOnePixelStream_s2mPipe_valid;
      end
      if(compareStage_counterOnePixelStream_valid) begin
        compareStage_counterOnePixelStream_rValid <= 1'b1;
      end
      if(compareStage_counterOnePixelStream_s2mPipe_ready) begin
        compareStage_counterOnePixelStream_rValid <= 1'b0;
      end
      if(compareStage_counterOnePixelStream_s2mPipe_ready) begin
        compareStage_counterOnePixelStream_s2mPipe_rValid <= compareStage_counterOnePixelStream_s2mPipe_valid;
      end
      if(compareStage_mainTwoPixelStream_valid) begin
        compareStage_mainTwoPixelStream_rValid <= 1'b1;
      end
      if(compareStage_mainTwoPixelStream_s2mPipe_ready) begin
        compareStage_mainTwoPixelStream_rValid <= 1'b0;
      end
      if(compareStage_mainTwoPixelStream_s2mPipe_ready) begin
        compareStage_mainTwoPixelStream_s2mPipe_rValid <= compareStage_mainTwoPixelStream_s2mPipe_valid;
      end
      if(compareStage_counterTwoPixelStream_valid) begin
        compareStage_counterTwoPixelStream_rValid <= 1'b1;
      end
      if(compareStage_counterTwoPixelStream_s2mPipe_ready) begin
        compareStage_counterTwoPixelStream_rValid <= 1'b0;
      end
      if(compareStage_counterTwoPixelStream_s2mPipe_ready) begin
        compareStage_counterTwoPixelStream_s2mPipe_rValid <= compareStage_counterTwoPixelStream_s2mPipe_valid;
      end
      if(compareStage_oddRowPixelStream_valid) begin
        compareStage_oddRowPixelStream_rValid <= 1'b1;
      end
      if(compareStage_oddRowPixelStream_s2mPipe_ready) begin
        compareStage_oddRowPixelStream_rValid <= 1'b0;
      end
      if(compareStage_oddRowPixelStream_s2mPipe_ready) begin
        compareStage_oddRowPixelStream_s2mPipe_rValid <= compareStage_oddRowPixelStream_s2mPipe_valid;
      end
      if(compareStage_controlPipe_translated_valid) begin
        compareStage_controlPipe_translated_rValid <= 1'b1;
      end
      if(compareStage_controlPipe_translated_s2mPipe_ready) begin
        compareStage_controlPipe_translated_rValid <= 1'b0;
      end
      if(compareStage_controlPipe_translated_s2mPipe_ready) begin
        compareStage_controlPipe_translated_s2mPipe_rValid <= compareStage_controlPipe_translated_s2mPipe_valid;
      end
      if(diffStage_mainOnePixelStream_valid) begin
        diffStage_mainOnePixelStream_rValid <= 1'b1;
      end
      if(diffStage_mainOnePixelStream_s2mPipe_ready) begin
        diffStage_mainOnePixelStream_rValid <= 1'b0;
      end
      if(diffStage_mainOnePixelStream_s2mPipe_ready) begin
        diffStage_mainOnePixelStream_s2mPipe_rValid <= diffStage_mainOnePixelStream_s2mPipe_valid;
      end
      if(diffStage_counterOnePixelStream_valid) begin
        diffStage_counterOnePixelStream_rValid <= 1'b1;
      end
      if(diffStage_counterOnePixelStream_s2mPipe_ready) begin
        diffStage_counterOnePixelStream_rValid <= 1'b0;
      end
      if(diffStage_counterOnePixelStream_s2mPipe_ready) begin
        diffStage_counterOnePixelStream_s2mPipe_rValid <= diffStage_counterOnePixelStream_s2mPipe_valid;
      end
      if(diffStage_mainTwoPixelStream_valid) begin
        diffStage_mainTwoPixelStream_rValid <= 1'b1;
      end
      if(diffStage_mainTwoPixelStream_s2mPipe_ready) begin
        diffStage_mainTwoPixelStream_rValid <= 1'b0;
      end
      if(diffStage_mainTwoPixelStream_s2mPipe_ready) begin
        diffStage_mainTwoPixelStream_s2mPipe_rValid <= diffStage_mainTwoPixelStream_s2mPipe_valid;
      end
      if(diffStage_counterTwoPixelStream_valid) begin
        diffStage_counterTwoPixelStream_rValid <= 1'b1;
      end
      if(diffStage_counterTwoPixelStream_s2mPipe_ready) begin
        diffStage_counterTwoPixelStream_rValid <= 1'b0;
      end
      if(diffStage_counterTwoPixelStream_s2mPipe_ready) begin
        diffStage_counterTwoPixelStream_s2mPipe_rValid <= diffStage_counterTwoPixelStream_s2mPipe_valid;
      end
      if(diffStage_oddRowPixelStream_valid) begin
        diffStage_oddRowPixelStream_rValid <= 1'b1;
      end
      if(diffStage_oddRowPixelStream_s2mPipe_ready) begin
        diffStage_oddRowPixelStream_rValid <= 1'b0;
      end
      if(diffStage_oddRowPixelStream_s2mPipe_ready) begin
        diffStage_oddRowPixelStream_s2mPipe_rValid <= diffStage_oddRowPixelStream_s2mPipe_valid;
      end
      if(diffStage_controlPipe_fork_io_outputs_0_translated_valid) begin
        diffStage_controlPipe_fork_io_outputs_0_translated_rValid <= 1'b1;
      end
      if(diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_ready) begin
        diffStage_controlPipe_fork_io_outputs_0_translated_rValid <= 1'b0;
      end
      if(diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_ready) begin
        diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rValid <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_valid;
      end
      if(resultStage_pixelStream_valid) begin
        resultStage_pixelStream_rValid <= 1'b1;
      end
      if(resultStage_pixelStream_s2mPipe_ready) begin
        resultStage_pixelStream_rValid <= 1'b0;
      end
      if(resultStage_pixelStream_s2mPipe_ready) begin
        resultStage_pixelStream_s2mPipe_rValid <= resultStage_pixelStream_s2mPipe_valid;
      end
      if(pixelsStream_valid) begin
        pixelsStream_rValid <= 1'b1;
      end
      if(pixelsStream_s2mPipe_ready) begin
        pixelsStream_rValid <= 1'b0;
      end
      if(pixelsStream_s2mPipe_ready) begin
        pixelsStream_s2mPipe_rValid <= pixelsStream_s2mPipe_valid;
      end
      if(when_SuperResolutionPart2_l761) begin
        if(when_SuperResolutionPart2_l763) begin
          outReachRowEnd <= 1'b1;
        end
        if(when_SuperResolutionPart2_l764) begin
          outReachFinalRow <= 1'b1;
        end
        if(when_SuperResolutionPart2_l766) begin
          if(outReachFinalRow) begin
            startRead <= 1'b0;
            readDone <= 1'b1;
            outReachRowEnd <= 1'b0;
            outReachFinalRow <= 1'b0;
          end else begin
            outReachRowEnd <= 1'b0;
          end
        end
        if(controlStream_fire_7) begin
          if(outReachRowEnd) begin
            outReachRowEnd <= 1'b0;
            if(when_SuperResolutionPart2_l783) begin
              oneInFourOutRow <= 1'b1;
            end else begin
              oneInFourOutRow <= 1'b0;
            end
            if(when_SuperResolutionPart2_l785) begin
              twoInFourOutRow <= 1'b1;
            end else begin
              twoInFourOutRow <= 1'b0;
            end
            if(when_SuperResolutionPart2_l787) begin
              threeInFourOutRow <= 1'b1;
            end else begin
              threeInFourOutRow <= 1'b0;
            end
            if(when_SuperResolutionPart2_l789) begin
              zeroInFourOutRow <= 1'b1;
            end else begin
              zeroInFourOutRow <= 1'b0;
            end
          end
          if(when_SuperResolutionPart2_l793) begin
            oneInFourOutPixelAddr <= 1'b1;
          end
          if(oneInFourOutPixelAddr) begin
            oneInFourOutPixelAddr <= 1'b0;
          end
          if(when_SuperResolutionPart2_l796) begin
            twoInFourOutPixelAddr <= 1'b1;
          end
          if(twoInFourOutPixelAddr) begin
            twoInFourOutPixelAddr <= 1'b0;
          end
          if(when_SuperResolutionPart2_l799) begin
            threeInFourOutPixelAddr <= 1'b1;
          end
          if(threeInFourOutPixelAddr) begin
            threeInFourOutPixelAddr <= 1'b0;
          end
          if(when_SuperResolutionPart2_l802) begin
            zeroInFourOutPixelAddr <= 1'b1;
          end
          if(zeroInFourOutPixelAddr) begin
            zeroInFourOutPixelAddr <= 1'b0;
          end
        end
      end
      controlStateMachine_stateReg <= controlStateMachine_stateNext;
      case(controlStateMachine_stateReg)
        controlStateMachine_enumDef_4_HOLD : begin
          if(zeroInFourOutRow) begin
            if(passPixels_fire_13) begin
              if(!threeInFourOutPixelAddr) begin
                holdWillPassToHoldCaseTwo <= 1'b1;
              end
            end
          end else begin
            if(!twoInFourOutRow) begin
              if(threeInFourOutRow) begin
                if(passPixels_fire_15) begin
                  if(threeInFourOutPixelAddr) begin
                    if(willHoldToTwice) begin
                      willHoldToTwice <= 1'b0;
                    end
                  end
                end
              end
            end
          end
          if(passPixels_fire_16) begin
            if(when_SuperResolutionPart2_l560) begin
              willHoldToTwice <= 1'b1;
            end else begin
              willHoldToTwice <= 1'b0;
            end
          end
        end
        controlStateMachine_enumDef_4_PASS : begin
          if(controlStream_fire_8) begin
            if(!oneInFourOutPixelAddr) begin
              if(twoInFourOutPixelAddr) begin
                if(oneInFourOutRow) begin
                  if(when_SuperResolutionPart2_l585) begin
                    willOnceToHoldCaseOne <= 1'b1;
                  end
                end else begin
                  if(twoInFourOutRow) begin
                    if(when_SuperResolutionPart2_l588) begin
                      willOnceToHoldCaseTwo <= 1'b1;
                    end
                  end else begin
                    if(when_SuperResolutionPart2_l590) begin
                      holdWillPassToHoldCaseTwo <= 1'b0;
                    end
                  end
                end
              end
            end
            willPassToHoldCaseOne <= 1'b0;
            willPassToHoldCaseTwo <= 1'b0;
          end
          if(when_SuperResolutionPart2_l602) begin
            willPassToHoldCaseOne <= 1'b1;
          end
          if(when_SuperResolutionPart2_l603) begin
            willPassToHoldCaseOne <= 1'b1;
          end
          if(when_SuperResolutionPart2_l605) begin
            willPassToHoldCaseTwo <= 1'b1;
          end
          if(when_SuperResolutionPart2_l606) begin
            willPassToHoldCaseTwo <= 1'b1;
          end
          if(when_SuperResolutionPart2_l630) begin
            frameStart <= 1'b0;
          end
        end
        controlStateMachine_enumDef_4_ONCE : begin
          if(controlStream_fire_10) begin
            willOnceToHoldCaseOne <= 1'b0;
            willOnceToHoldCaseTwo <= 1'b0;
            willOnceToHoldCaseThree <= 1'b0;
          end
          if(when_SuperResolutionPart2_l662) begin
            willOnceToHoldCaseOne <= 1'b0;
            willOnceToHoldCaseTwo <= 1'b0;
          end
          if(when_SuperResolutionPart2_l667) begin
            willOnceToHoldCaseThree <= 1'b1;
          end
          if(when_SuperResolutionPart2_l668) begin
            willOnceToHoldCaseThree <= 1'b1;
          end
        end
        controlStateMachine_enumDef_4_TWICE : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(posedge clk) begin
    startIn_regNext <= startIn;
    startIn_regNext_1 <= startIn;
    startIn_regNext_2 <= startIn;
    startIn_regNext_3 <= startIn;
    startIn_regNext_4 <= startIn;
    startIn_regNext_5 <= startIn;
    startIn_regNext_6 <= startIn;
    startIn_regNext_7 <= startIn;
    startIn_regNext_8 <= startIn;
    startIn_regNext_9 <= startIn;
    startIn_regNext_10 <= startIn;
    startIn_regNext_11 <= startIn;
    startIn_regNext_12 <= startIn;
    startIn_regNext_13 <= startIn;
    startIn_regNext_14 <= startIn;
    startIn_regNext_15 <= startIn;
    startIn_regNext_16 <= startIn;
    if(pixelsIn_ready) begin
      pixelsIn_rData_pixel <= pixelsIn_payload_pixel;
      pixelsIn_rData_frameStart <= pixelsIn_payload_frameStart;
      pixelsIn_rData_rowEnd <= pixelsIn_payload_rowEnd;
    end
    if(pixelsIn_s2mPipe_ready) begin
      pixelsIn_s2mPipe_rData_pixel <= pixelsIn_s2mPipe_payload_pixel;
      pixelsIn_s2mPipe_rData_frameStart <= pixelsIn_s2mPipe_payload_frameStart;
      pixelsIn_s2mPipe_rData_rowEnd <= pixelsIn_s2mPipe_payload_rowEnd;
    end
    if(mainAddrOneStream_ready) begin
      mainAddrOneStream_rData <= mainAddrOneStream_payload;
    end
    if(mainAddrOneStream_s2mPipe_ready) begin
      mainAddrOneStream_s2mPipe_rData <= mainAddrOneStream_s2mPipe_payload;
    end
    if(CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_mainOnePixelStream_payload_1 <= CICC1851_readStage_mainOnePixelStream_payload;
    end
    if(CICC1851_1) begin
      CICC1851_readStage_mainOnePixelStream_payload_2 <= (CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_mainOnePixelStream_payload_1 : CICC1851_readStage_mainOnePixelStream_payload);
    end
    if(counterAddrOneStream_ready) begin
      counterAddrOneStream_rData <= counterAddrOneStream_payload;
    end
    if(counterAddrOneStream_s2mPipe_ready) begin
      counterAddrOneStream_s2mPipe_rData <= counterAddrOneStream_s2mPipe_payload;
    end
    if(CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_counterOnePixelStream_payload_1 <= CICC1851_readStage_counterOnePixelStream_payload;
    end
    if(CICC1851_2) begin
      CICC1851_readStage_counterOnePixelStream_payload_2 <= (CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_counterOnePixelStream_payload_1 : CICC1851_readStage_counterOnePixelStream_payload);
    end
    if(mainAddrTwoStream_ready) begin
      mainAddrTwoStream_rData <= mainAddrTwoStream_payload;
    end
    if(mainAddrTwoStream_s2mPipe_ready) begin
      mainAddrTwoStream_s2mPipe_rData <= mainAddrTwoStream_s2mPipe_payload;
    end
    if(CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_mainTwoPixelStream_payload_1 <= CICC1851_readStage_mainTwoPixelStream_payload;
    end
    if(CICC1851_3) begin
      CICC1851_readStage_mainTwoPixelStream_payload_2 <= (CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_mainTwoPixelStream_payload_1 : CICC1851_readStage_mainTwoPixelStream_payload);
    end
    if(counterAddrTwoStream_ready) begin
      counterAddrTwoStream_rData <= counterAddrTwoStream_payload;
    end
    if(counterAddrTwoStream_s2mPipe_ready) begin
      counterAddrTwoStream_s2mPipe_rData <= counterAddrTwoStream_s2mPipe_payload;
    end
    if(CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_counterTwoPixelStream_payload_1 <= CICC1851_readStage_counterTwoPixelStream_payload;
    end
    if(CICC1851_4) begin
      CICC1851_readStage_counterTwoPixelStream_payload_2 <= (CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_counterTwoPixelStream_payload_1 : CICC1851_readStage_counterTwoPixelStream_payload);
    end
    if(oddAddrStream_ready) begin
      oddAddrStream_rData <= oddAddrStream_payload;
    end
    if(oddAddrStream_s2mPipe_ready) begin
      oddAddrStream_s2mPipe_rData <= oddAddrStream_s2mPipe_payload;
    end
    if(CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_oddRowPixelStream_payload_1 <= CICC1851_readStage_oddRowPixelStream_payload;
    end
    if(CICC1851_5) begin
      CICC1851_readStage_oddRowPixelStream_payload_2 <= (CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_oddRowPixelStream_payload_1 : CICC1851_readStage_oddRowPixelStream_payload);
    end
    if(controlStream_ready) begin
      controlStream_rData_frameStart <= controlStream_payload_frameStart;
      controlStream_rData_rowEnd <= controlStream_payload_rowEnd;
      controlStream_rData_passMode <= controlStream_payload_passMode;
      controlStream_rData_passValid <= controlStream_payload_passValid;
      controlStream_rData_onceMode <= controlStream_payload_onceMode;
      controlStream_rData_onceValid <= controlStream_payload_onceValid;
      controlStream_rData_mainCompare <= controlStream_payload_mainCompare;
      controlStream_rData_counterCompare <= controlStream_payload_counterCompare;
      controlStream_rData_mainDiff <= controlStream_payload_mainDiff;
      controlStream_rData_counterDiff <= controlStream_payload_counterDiff;
      controlStream_rData_twiceCompValid <= controlStream_payload_twiceCompValid;
      controlStream_rData_twiceMode <= controlStream_payload_twiceMode;
      controlStream_rData_inpValidFlag <= controlStream_payload_inpValidFlag;
      controlStream_rData_oddValid <= controlStream_payload_oddValid;
    end
    if(controlStream_s2mPipe_ready) begin
      controlStream_s2mPipe_rData_frameStart <= controlStream_s2mPipe_payload_frameStart;
      controlStream_s2mPipe_rData_rowEnd <= controlStream_s2mPipe_payload_rowEnd;
      controlStream_s2mPipe_rData_passMode <= controlStream_s2mPipe_payload_passMode;
      controlStream_s2mPipe_rData_passValid <= controlStream_s2mPipe_payload_passValid;
      controlStream_s2mPipe_rData_onceMode <= controlStream_s2mPipe_payload_onceMode;
      controlStream_s2mPipe_rData_onceValid <= controlStream_s2mPipe_payload_onceValid;
      controlStream_s2mPipe_rData_mainCompare <= controlStream_s2mPipe_payload_mainCompare;
      controlStream_s2mPipe_rData_counterCompare <= controlStream_s2mPipe_payload_counterCompare;
      controlStream_s2mPipe_rData_mainDiff <= controlStream_s2mPipe_payload_mainDiff;
      controlStream_s2mPipe_rData_counterDiff <= controlStream_s2mPipe_payload_counterDiff;
      controlStream_s2mPipe_rData_twiceCompValid <= controlStream_s2mPipe_payload_twiceCompValid;
      controlStream_s2mPipe_rData_twiceMode <= controlStream_s2mPipe_payload_twiceMode;
      controlStream_s2mPipe_rData_inpValidFlag <= controlStream_s2mPipe_payload_inpValidFlag;
      controlStream_s2mPipe_rData_oddValid <= controlStream_s2mPipe_payload_oddValid;
    end
    if(controlStream_s2mPipe_m2sPipe_ready) begin
      controlStream_s2mPipe_m2sPipe_rData_frameStart <= controlStream_s2mPipe_m2sPipe_payload_frameStart;
      controlStream_s2mPipe_m2sPipe_rData_rowEnd <= controlStream_s2mPipe_m2sPipe_payload_rowEnd;
      controlStream_s2mPipe_m2sPipe_rData_passMode <= controlStream_s2mPipe_m2sPipe_payload_passMode;
      controlStream_s2mPipe_m2sPipe_rData_passValid <= controlStream_s2mPipe_m2sPipe_payload_passValid;
      controlStream_s2mPipe_m2sPipe_rData_onceMode <= controlStream_s2mPipe_m2sPipe_payload_onceMode;
      controlStream_s2mPipe_m2sPipe_rData_onceValid <= controlStream_s2mPipe_m2sPipe_payload_onceValid;
      controlStream_s2mPipe_m2sPipe_rData_mainCompare <= controlStream_s2mPipe_m2sPipe_payload_mainCompare;
      controlStream_s2mPipe_m2sPipe_rData_counterCompare <= controlStream_s2mPipe_m2sPipe_payload_counterCompare;
      controlStream_s2mPipe_m2sPipe_rData_mainDiff <= controlStream_s2mPipe_m2sPipe_payload_mainDiff;
      controlStream_s2mPipe_m2sPipe_rData_counterDiff <= controlStream_s2mPipe_m2sPipe_payload_counterDiff;
      controlStream_s2mPipe_m2sPipe_rData_twiceCompValid <= controlStream_s2mPipe_m2sPipe_payload_twiceCompValid;
      controlStream_s2mPipe_m2sPipe_rData_twiceMode <= controlStream_s2mPipe_m2sPipe_payload_twiceMode;
      controlStream_s2mPipe_m2sPipe_rData_inpValidFlag <= controlStream_s2mPipe_m2sPipe_payload_inpValidFlag;
      controlStream_s2mPipe_m2sPipe_rData_oddValid <= controlStream_s2mPipe_m2sPipe_payload_oddValid;
    end
    if(controlStream_s2mPipe_m2sPipe_m2sPipe_ready) begin
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_frameStart <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_frameStart;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_rowEnd <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_rowEnd;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_passMode <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passMode;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_passValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_onceMode <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceMode;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_onceValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_twiceCompValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceCompValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_twiceMode <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceMode;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_inpValidFlag <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_inpValidFlag;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_oddValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_oddValid;
    end
    if(controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready) begin
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_frameStart <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_frameStart;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_rowEnd <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_rowEnd;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_passMode <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_passMode;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_passValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_passValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_onceMode <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_onceMode;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_onceValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_onceValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_twiceCompValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_twiceCompValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_twiceMode <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_twiceMode;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_inpValidFlag <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_inpValidFlag;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_oddValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_oddValid;
    end
    if(readStage_mainOnePixelStream_ready) begin
      readStage_mainOnePixelStream_rData <= readStage_mainOnePixelStream_payload;
    end
    if(readStage_mainOnePixelStream_s2mPipe_ready) begin
      readStage_mainOnePixelStream_s2mPipe_rData <= readStage_mainOnePixelStream_s2mPipe_payload;
    end
    if(readStage_counterOnePixelStream_ready) begin
      readStage_counterOnePixelStream_rData <= readStage_counterOnePixelStream_payload;
    end
    if(readStage_counterOnePixelStream_s2mPipe_ready) begin
      readStage_counterOnePixelStream_s2mPipe_rData <= readStage_counterOnePixelStream_s2mPipe_payload;
    end
    if(readStage_mainTwoPixelStream_ready) begin
      readStage_mainTwoPixelStream_rData <= readStage_mainTwoPixelStream_payload;
    end
    if(readStage_mainTwoPixelStream_s2mPipe_ready) begin
      readStage_mainTwoPixelStream_s2mPipe_rData <= readStage_mainTwoPixelStream_s2mPipe_payload;
    end
    if(readStage_counterTwoPixelStream_ready) begin
      readStage_counterTwoPixelStream_rData <= readStage_counterTwoPixelStream_payload;
    end
    if(readStage_counterTwoPixelStream_s2mPipe_ready) begin
      readStage_counterTwoPixelStream_s2mPipe_rData <= readStage_counterTwoPixelStream_s2mPipe_payload;
    end
    if(readStage_oddRowPixelStream_ready) begin
      readStage_oddRowPixelStream_rData <= readStage_oddRowPixelStream_payload;
    end
    if(readStage_oddRowPixelStream_s2mPipe_ready) begin
      readStage_oddRowPixelStream_s2mPipe_rData <= readStage_oddRowPixelStream_s2mPipe_payload;
    end
    if(readStage_controlPipe_translated_ready) begin
      readStage_controlPipe_translated_rData_frameStart <= readStage_controlPipe_translated_payload_frameStart;
      readStage_controlPipe_translated_rData_rowEnd <= readStage_controlPipe_translated_payload_rowEnd;
      readStage_controlPipe_translated_rData_passMode <= readStage_controlPipe_translated_payload_passMode;
      readStage_controlPipe_translated_rData_passValid <= readStage_controlPipe_translated_payload_passValid;
      readStage_controlPipe_translated_rData_onceMode <= readStage_controlPipe_translated_payload_onceMode;
      readStage_controlPipe_translated_rData_onceValid <= readStage_controlPipe_translated_payload_onceValid;
      readStage_controlPipe_translated_rData_mainCompare <= readStage_controlPipe_translated_payload_mainCompare;
      readStage_controlPipe_translated_rData_counterCompare <= readStage_controlPipe_translated_payload_counterCompare;
      readStage_controlPipe_translated_rData_mainDiff <= readStage_controlPipe_translated_payload_mainDiff;
      readStage_controlPipe_translated_rData_counterDiff <= readStage_controlPipe_translated_payload_counterDiff;
      readStage_controlPipe_translated_rData_twiceCompValid <= readStage_controlPipe_translated_payload_twiceCompValid;
      readStage_controlPipe_translated_rData_twiceMode <= readStage_controlPipe_translated_payload_twiceMode;
      readStage_controlPipe_translated_rData_inpValidFlag <= readStage_controlPipe_translated_payload_inpValidFlag;
      readStage_controlPipe_translated_rData_oddValid <= readStage_controlPipe_translated_payload_oddValid;
    end
    if(readStage_controlPipe_translated_s2mPipe_ready) begin
      readStage_controlPipe_translated_s2mPipe_rData_frameStart <= readStage_controlPipe_translated_s2mPipe_payload_frameStart;
      readStage_controlPipe_translated_s2mPipe_rData_rowEnd <= readStage_controlPipe_translated_s2mPipe_payload_rowEnd;
      readStage_controlPipe_translated_s2mPipe_rData_passMode <= readStage_controlPipe_translated_s2mPipe_payload_passMode;
      readStage_controlPipe_translated_s2mPipe_rData_passValid <= readStage_controlPipe_translated_s2mPipe_payload_passValid;
      readStage_controlPipe_translated_s2mPipe_rData_onceMode <= readStage_controlPipe_translated_s2mPipe_payload_onceMode;
      readStage_controlPipe_translated_s2mPipe_rData_onceValid <= readStage_controlPipe_translated_s2mPipe_payload_onceValid;
      readStage_controlPipe_translated_s2mPipe_rData_mainCompare <= readStage_controlPipe_translated_s2mPipe_payload_mainCompare;
      readStage_controlPipe_translated_s2mPipe_rData_counterCompare <= readStage_controlPipe_translated_s2mPipe_payload_counterCompare;
      readStage_controlPipe_translated_s2mPipe_rData_mainDiff <= readStage_controlPipe_translated_s2mPipe_payload_mainDiff;
      readStage_controlPipe_translated_s2mPipe_rData_counterDiff <= readStage_controlPipe_translated_s2mPipe_payload_counterDiff;
      readStage_controlPipe_translated_s2mPipe_rData_twiceCompValid <= readStage_controlPipe_translated_s2mPipe_payload_twiceCompValid;
      readStage_controlPipe_translated_s2mPipe_rData_twiceMode <= readStage_controlPipe_translated_s2mPipe_payload_twiceMode;
      readStage_controlPipe_translated_s2mPipe_rData_inpValidFlag <= readStage_controlPipe_translated_s2mPipe_payload_inpValidFlag;
      readStage_controlPipe_translated_s2mPipe_rData_oddValid <= readStage_controlPipe_translated_s2mPipe_payload_oddValid;
    end
    if(compareStage_mainOnePixelStream_ready) begin
      compareStage_mainOnePixelStream_rData <= compareStage_mainOnePixelStream_payload;
    end
    if(compareStage_mainOnePixelStream_s2mPipe_ready) begin
      compareStage_mainOnePixelStream_s2mPipe_rData <= compareStage_mainOnePixelStream_s2mPipe_payload;
    end
    if(compareStage_counterOnePixelStream_ready) begin
      compareStage_counterOnePixelStream_rData <= compareStage_counterOnePixelStream_payload;
    end
    if(compareStage_counterOnePixelStream_s2mPipe_ready) begin
      compareStage_counterOnePixelStream_s2mPipe_rData <= compareStage_counterOnePixelStream_s2mPipe_payload;
    end
    if(compareStage_mainTwoPixelStream_ready) begin
      compareStage_mainTwoPixelStream_rData <= compareStage_mainTwoPixelStream_payload;
    end
    if(compareStage_mainTwoPixelStream_s2mPipe_ready) begin
      compareStage_mainTwoPixelStream_s2mPipe_rData <= compareStage_mainTwoPixelStream_s2mPipe_payload;
    end
    if(compareStage_counterTwoPixelStream_ready) begin
      compareStage_counterTwoPixelStream_rData <= compareStage_counterTwoPixelStream_payload;
    end
    if(compareStage_counterTwoPixelStream_s2mPipe_ready) begin
      compareStage_counterTwoPixelStream_s2mPipe_rData <= compareStage_counterTwoPixelStream_s2mPipe_payload;
    end
    if(compareStage_oddRowPixelStream_ready) begin
      compareStage_oddRowPixelStream_rData <= compareStage_oddRowPixelStream_payload;
    end
    if(compareStage_oddRowPixelStream_s2mPipe_ready) begin
      compareStage_oddRowPixelStream_s2mPipe_rData <= compareStage_oddRowPixelStream_s2mPipe_payload;
    end
    if(compareStage_controlPipe_translated_ready) begin
      compareStage_controlPipe_translated_rData_frameStart <= compareStage_controlPipe_translated_payload_frameStart;
      compareStage_controlPipe_translated_rData_rowEnd <= compareStage_controlPipe_translated_payload_rowEnd;
      compareStage_controlPipe_translated_rData_passMode <= compareStage_controlPipe_translated_payload_passMode;
      compareStage_controlPipe_translated_rData_passValid <= compareStage_controlPipe_translated_payload_passValid;
      compareStage_controlPipe_translated_rData_onceMode <= compareStage_controlPipe_translated_payload_onceMode;
      compareStage_controlPipe_translated_rData_onceValid <= compareStage_controlPipe_translated_payload_onceValid;
      compareStage_controlPipe_translated_rData_mainCompare <= compareStage_controlPipe_translated_payload_mainCompare;
      compareStage_controlPipe_translated_rData_counterCompare <= compareStage_controlPipe_translated_payload_counterCompare;
      compareStage_controlPipe_translated_rData_mainDiff <= compareStage_controlPipe_translated_payload_mainDiff;
      compareStage_controlPipe_translated_rData_counterDiff <= compareStage_controlPipe_translated_payload_counterDiff;
      compareStage_controlPipe_translated_rData_twiceCompValid <= compareStage_controlPipe_translated_payload_twiceCompValid;
      compareStage_controlPipe_translated_rData_twiceMode <= compareStage_controlPipe_translated_payload_twiceMode;
      compareStage_controlPipe_translated_rData_inpValidFlag <= compareStage_controlPipe_translated_payload_inpValidFlag;
      compareStage_controlPipe_translated_rData_oddValid <= compareStage_controlPipe_translated_payload_oddValid;
    end
    if(compareStage_controlPipe_translated_s2mPipe_ready) begin
      compareStage_controlPipe_translated_s2mPipe_rData_frameStart <= compareStage_controlPipe_translated_s2mPipe_payload_frameStart;
      compareStage_controlPipe_translated_s2mPipe_rData_rowEnd <= compareStage_controlPipe_translated_s2mPipe_payload_rowEnd;
      compareStage_controlPipe_translated_s2mPipe_rData_passMode <= compareStage_controlPipe_translated_s2mPipe_payload_passMode;
      compareStage_controlPipe_translated_s2mPipe_rData_passValid <= compareStage_controlPipe_translated_s2mPipe_payload_passValid;
      compareStage_controlPipe_translated_s2mPipe_rData_onceMode <= compareStage_controlPipe_translated_s2mPipe_payload_onceMode;
      compareStage_controlPipe_translated_s2mPipe_rData_onceValid <= compareStage_controlPipe_translated_s2mPipe_payload_onceValid;
      compareStage_controlPipe_translated_s2mPipe_rData_mainCompare <= compareStage_controlPipe_translated_s2mPipe_payload_mainCompare;
      compareStage_controlPipe_translated_s2mPipe_rData_counterCompare <= compareStage_controlPipe_translated_s2mPipe_payload_counterCompare;
      compareStage_controlPipe_translated_s2mPipe_rData_mainDiff <= compareStage_controlPipe_translated_s2mPipe_payload_mainDiff;
      compareStage_controlPipe_translated_s2mPipe_rData_counterDiff <= compareStage_controlPipe_translated_s2mPipe_payload_counterDiff;
      compareStage_controlPipe_translated_s2mPipe_rData_twiceCompValid <= compareStage_controlPipe_translated_s2mPipe_payload_twiceCompValid;
      compareStage_controlPipe_translated_s2mPipe_rData_twiceMode <= compareStage_controlPipe_translated_s2mPipe_payload_twiceMode;
      compareStage_controlPipe_translated_s2mPipe_rData_inpValidFlag <= compareStage_controlPipe_translated_s2mPipe_payload_inpValidFlag;
      compareStage_controlPipe_translated_s2mPipe_rData_oddValid <= compareStage_controlPipe_translated_s2mPipe_payload_oddValid;
    end
    if(diffStage_mainOnePixelStream_ready) begin
      diffStage_mainOnePixelStream_rData <= diffStage_mainOnePixelStream_payload;
    end
    if(diffStage_mainOnePixelStream_s2mPipe_ready) begin
      diffStage_mainOnePixelStream_s2mPipe_rData <= diffStage_mainOnePixelStream_s2mPipe_payload;
    end
    if(diffStage_counterOnePixelStream_ready) begin
      diffStage_counterOnePixelStream_rData <= diffStage_counterOnePixelStream_payload;
    end
    if(diffStage_counterOnePixelStream_s2mPipe_ready) begin
      diffStage_counterOnePixelStream_s2mPipe_rData <= diffStage_counterOnePixelStream_s2mPipe_payload;
    end
    if(diffStage_mainTwoPixelStream_ready) begin
      diffStage_mainTwoPixelStream_rData <= diffStage_mainTwoPixelStream_payload;
    end
    if(diffStage_mainTwoPixelStream_s2mPipe_ready) begin
      diffStage_mainTwoPixelStream_s2mPipe_rData <= diffStage_mainTwoPixelStream_s2mPipe_payload;
    end
    if(diffStage_counterTwoPixelStream_ready) begin
      diffStage_counterTwoPixelStream_rData <= diffStage_counterTwoPixelStream_payload;
    end
    if(diffStage_counterTwoPixelStream_s2mPipe_ready) begin
      diffStage_counterTwoPixelStream_s2mPipe_rData <= diffStage_counterTwoPixelStream_s2mPipe_payload;
    end
    if(diffStage_oddRowPixelStream_ready) begin
      diffStage_oddRowPixelStream_rData <= diffStage_oddRowPixelStream_payload;
    end
    if(diffStage_oddRowPixelStream_s2mPipe_ready) begin
      diffStage_oddRowPixelStream_s2mPipe_rData <= diffStage_oddRowPixelStream_s2mPipe_payload;
    end
    if(diffStage_controlPipe_fork_io_outputs_0_translated_ready) begin
      diffStage_controlPipe_fork_io_outputs_0_translated_rData_frameStart <= diffStage_controlPipe_fork_io_outputs_0_translated_payload_frameStart;
      diffStage_controlPipe_fork_io_outputs_0_translated_rData_rowEnd <= diffStage_controlPipe_fork_io_outputs_0_translated_payload_rowEnd;
      diffStage_controlPipe_fork_io_outputs_0_translated_rData_passMode <= diffStage_controlPipe_fork_io_outputs_0_translated_payload_passMode;
      diffStage_controlPipe_fork_io_outputs_0_translated_rData_passValid <= diffStage_controlPipe_fork_io_outputs_0_translated_payload_passValid;
      diffStage_controlPipe_fork_io_outputs_0_translated_rData_onceMode <= diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceMode;
      diffStage_controlPipe_fork_io_outputs_0_translated_rData_onceValid <= diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceValid;
      diffStage_controlPipe_fork_io_outputs_0_translated_rData_mainCompare <= diffStage_controlPipe_fork_io_outputs_0_translated_payload_mainCompare;
      diffStage_controlPipe_fork_io_outputs_0_translated_rData_counterCompare <= diffStage_controlPipe_fork_io_outputs_0_translated_payload_counterCompare;
      diffStage_controlPipe_fork_io_outputs_0_translated_rData_mainDiff <= diffStage_controlPipe_fork_io_outputs_0_translated_payload_mainDiff;
      diffStage_controlPipe_fork_io_outputs_0_translated_rData_counterDiff <= diffStage_controlPipe_fork_io_outputs_0_translated_payload_counterDiff;
      diffStage_controlPipe_fork_io_outputs_0_translated_rData_twiceCompValid <= diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceCompValid;
      diffStage_controlPipe_fork_io_outputs_0_translated_rData_twiceMode <= diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceMode;
      diffStage_controlPipe_fork_io_outputs_0_translated_rData_inpValidFlag <= diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag;
      diffStage_controlPipe_fork_io_outputs_0_translated_rData_oddValid <= diffStage_controlPipe_fork_io_outputs_0_translated_payload_oddValid;
    end
    if(diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_ready) begin
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_frameStart <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_frameStart;
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_rowEnd <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_rowEnd;
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_passMode <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_passMode;
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_passValid <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_passValid;
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_onceMode <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_onceMode;
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_onceValid <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_onceValid;
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_mainCompare <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_mainCompare;
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_counterCompare <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_counterCompare;
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_mainDiff <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_mainDiff;
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_counterDiff <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_counterDiff;
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_twiceCompValid <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_twiceCompValid;
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_twiceMode <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_twiceMode;
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_inpValidFlag <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_inpValidFlag;
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_oddValid <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_oddValid;
    end
    if(resultStage_pixelStream_ready) begin
      resultStage_pixelStream_rData <= resultStage_pixelStream_payload;
    end
    if(resultStage_pixelStream_s2mPipe_ready) begin
      resultStage_pixelStream_s2mPipe_rData <= resultStage_pixelStream_s2mPipe_payload;
    end
    if(pixelsStream_ready) begin
      pixelsStream_rData_pixel <= pixelsStream_payload_pixel;
      pixelsStream_rData_frameStart <= pixelsStream_payload_frameStart;
      pixelsStream_rData_rowEnd <= pixelsStream_payload_rowEnd;
      pixelsStream_rData_inpValid <= pixelsStream_payload_inpValid;
    end
    if(pixelsStream_s2mPipe_ready) begin
      pixelsStream_s2mPipe_rData_pixel <= pixelsStream_s2mPipe_payload_pixel;
      pixelsStream_s2mPipe_rData_frameStart <= pixelsStream_s2mPipe_payload_frameStart;
      pixelsStream_s2mPipe_rData_rowEnd <= pixelsStream_s2mPipe_payload_rowEnd;
      pixelsStream_s2mPipe_rData_inpValid <= pixelsStream_s2mPipe_payload_inpValid;
    end
  end


endmodule

module SuperResolutionPart1_1 (
  input               pixelsIn_valid,
  output reg          pixelsIn_ready,
  input      [7:0]    pixelsIn_payload_pixel,
  input               pixelsIn_payload_frameStart,
  input               pixelsIn_payload_rowEnd,
  input               startIn,
  input               inpTwoDoneIn,
  input               inpThreeDoneIn,
  output reg          pixelsOut_valid,
  input               pixelsOut_ready,
  output reg [7:0]    pixelsOut_payload_pixel,
  output reg          pixelsOut_payload_frameStart,
  output reg          pixelsOut_payload_rowEnd,
  output reg          startOut,
  output reg          inpDoneOut,
  input      [7:0]    thresholdIn,
  input      [9:0]    widthIn,
  input      [9:0]    heightIn,
  input               clk,
  input               resetn
);
  localparam controlStateMachine_enumDef_3_BOOT = 3'd0;
  localparam controlStateMachine_enumDef_3_HOLD = 3'd1;
  localparam controlStateMachine_enumDef_3_PASS = 3'd2;
  localparam controlStateMachine_enumDef_3_ONCE = 3'd3;
  localparam controlStateMachine_enumDef_3_TWICE = 3'd4;

  wire                diffStage_controlPipe_fork_io_outputs_0_ready;
  reg        [7:0]    CICC1851_lineBufferOne_port0;
  reg        [7:0]    CICC1851_lineBufferOne_port1;
  reg        [7:0]    CICC1851_lineBufferTwo_port0;
  reg        [7:0]    CICC1851_lineBufferTwo_port1;
  wire                diffStage_controlPipe_fork_io_input_ready;
  wire                diffStage_controlPipe_fork_io_outputs_0_valid;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_frameStart;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_rowEnd;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_passMode;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_passValid;
  wire       [2:0]    diffStage_controlPipe_fork_io_outputs_0_payload_onceMode;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_onceValid;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_mainCompare;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_counterCompare;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_payload_mainDiff;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_payload_counterDiff;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_twiceCompValid;
  wire       [2:0]    diffStage_controlPipe_fork_io_outputs_0_payload_twiceMode;
  wire                diffStage_controlPipe_fork_io_outputs_1_valid;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_frameStart;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_rowEnd;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_passMode;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_passValid;
  wire       [2:0]    diffStage_controlPipe_fork_io_outputs_1_payload_onceMode;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_onceValid;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_mainCompare;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_counterCompare;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_twiceCompValid;
  wire       [2:0]    diffStage_controlPipe_fork_io_outputs_1_payload_twiceMode;
  wire       [9:0]    CICC1851_bufferRowCount_valueNext;
  wire       [0:0]    CICC1851_bufferRowCount_valueNext_1;
  wire       [9:0]    CICC1851_bufferWAddr_valueNext;
  wire       [0:0]    CICC1851_bufferWAddr_valueNext_1;
  wire       [10:0]   CICC1851_outPixelAddr_valueNext;
  wire       [0:0]    CICC1851_outPixelAddr_valueNext_1;
  wire       [10:0]   CICC1851_outRowCount_valueNext;
  wire       [0:0]    CICC1851_outRowCount_valueNext_1;
  wire       [10:0]   CICC1851_mainAddrOne;
  wire       [10:0]   CICC1851_counterAddrOne;
  wire       [10:0]   CICC1851_mainAddrTwo;
  wire       [10:0]   CICC1851_counterAddrTwo;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_1;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_2;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_3;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_4;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_5;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_6;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_7;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_8;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_9;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_10;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_11;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_12;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_13;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_14;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_15;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_16;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_17;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_18;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_19;
  wire       [9:0]    CICC1851_when_SuperResolutionPart1_l421;
  wire       [9:0]    CICC1851_when_SuperResolutionPart1_l422;
  wire       [10:0]   CICC1851_when_SuperResolutionPart1_l447;
  wire       [7:0]    CICC1851_lineBufferTwo_port;
  wire                CICC1851_lineBufferTwo_port_1;
  wire       [7:0]    CICC1851_lineBufferOne_port;
  wire                CICC1851_lineBufferOne_port_1;
  wire       [10:0]   CICC1851_when_SuperResolutionPart1_l482;
  wire       [10:0]   CICC1851_when_SuperResolutionPart1_l484;
  wire       [10:0]   CICC1851_when_SuperResolutionPart1_l489;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l498;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l498_1;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l500;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l500_1;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l500_2;
  wire       [2:0]    CICC1851_when_SuperResolutionPart1_l500_3;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l510;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l510_1;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l510_2;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l511;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l511_1;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l511_2;
  wire       [10:0]   CICC1851_when_SuperResolutionPart1_l537;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l542;
  wire       [10:0]   CICC1851_when_SuperResolutionPart1_l542_1;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l542_2;
  wire       [10:0]   CICC1851_mainAddrOne_1;
  wire       [10:0]   CICC1851_mainAddrOne_2;
  wire       [10:0]   CICC1851_counterAddrOne_1;
  wire       [10:0]   CICC1851_counterAddrOne_2;
  wire       [11:0]   CICC1851_counterAddrOne_3;
  wire       [11:0]   CICC1851_counterAddrOne_4;
  wire       [11:0]   CICC1851_counterAddrOne_5;
  wire       [1:0]    CICC1851_counterAddrOne_6;
  wire       [0:0]    CICC1851_controls_onceMode;
  wire       [10:0]   CICC1851_mainAddrTwo_1;
  wire       [10:0]   CICC1851_mainAddrTwo_2;
  wire       [10:0]   CICC1851_counterAddrTwo_1;
  wire       [10:0]   CICC1851_counterAddrTwo_2;
  wire       [11:0]   CICC1851_counterAddrTwo_3;
  wire       [11:0]   CICC1851_counterAddrTwo_4;
  wire       [11:0]   CICC1851_counterAddrTwo_5;
  wire       [1:0]    CICC1851_counterAddrTwo_6;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l563;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l563_1;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l563_2;
  wire       [2:0]    CICC1851_when_SuperResolutionPart1_l563_3;
  wire       [1:0]    CICC1851_controls_onceMode_1;
  wire       [1:0]    CICC1851_controls_onceMode_2;
  wire       [10:0]   CICC1851_mainAddrOne_3;
  wire       [10:0]   CICC1851_mainAddrTwo_3;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l578;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l578_1;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l578_2;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l579;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l579_1;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l579_2;
  wire       [10:0]   CICC1851_mainAddrOne_4;
  wire       [10:0]   CICC1851_mainAddrOne_5;
  wire       [10:0]   CICC1851_mainAddrOne_6;
  wire       [10:0]   CICC1851_mainAddrOne_7;
  wire       [11:0]   CICC1851_counterAddrOne_7;
  wire       [11:0]   CICC1851_counterAddrOne_8;
  wire       [11:0]   CICC1851_counterAddrOne_9;
  wire       [1:0]    CICC1851_counterAddrOne_10;
  wire       [10:0]   CICC1851_mainAddrTwo_4;
  wire       [10:0]   CICC1851_mainAddrTwo_5;
  wire       [10:0]   CICC1851_mainAddrTwo_6;
  wire       [10:0]   CICC1851_mainAddrTwo_7;
  wire       [11:0]   CICC1851_counterAddrTwo_7;
  wire       [11:0]   CICC1851_counterAddrTwo_8;
  wire       [11:0]   CICC1851_counterAddrTwo_9;
  wire       [1:0]    CICC1851_counterAddrTwo_10;
  wire       [10:0]   CICC1851_mainAddrOne_8;
  wire       [10:0]   CICC1851_mainAddrOne_9;
  wire       [10:0]   CICC1851_counterAddrTwo_11;
  wire       [10:0]   CICC1851_counterAddrTwo_12;
  wire       [10:0]   CICC1851_mainAddrTwo_8;
  wire       [10:0]   CICC1851_mainAddrTwo_9;
  wire       [10:0]   CICC1851_counterAddrOne_11;
  wire       [10:0]   CICC1851_counterAddrOne_12;
  wire       [11:0]   CICC1851_mainAddrTwo_10;
  wire       [11:0]   CICC1851_mainAddrTwo_11;
  wire       [11:0]   CICC1851_mainAddrTwo_12;
  wire       [1:0]    CICC1851_mainAddrTwo_13;
  wire       [11:0]   CICC1851_counterAddrOne_13;
  wire       [11:0]   CICC1851_counterAddrOne_14;
  wire       [11:0]   CICC1851_counterAddrOne_15;
  wire       [1:0]    CICC1851_counterAddrOne_16;
  wire       [10:0]   CICC1851_mainAddrTwo_14;
  wire       [10:0]   CICC1851_mainAddrTwo_15;
  wire       [10:0]   CICC1851_counterAddrOne_17;
  wire       [10:0]   CICC1851_counterAddrOne_18;
  wire       [10:0]   CICC1851_mainAddrOne_10;
  wire       [10:0]   CICC1851_mainAddrOne_11;
  wire       [10:0]   CICC1851_counterAddrTwo_13;
  wire       [10:0]   CICC1851_counterAddrTwo_14;
  wire       [11:0]   CICC1851_mainAddrOne_12;
  wire       [11:0]   CICC1851_mainAddrOne_13;
  wire       [11:0]   CICC1851_mainAddrOne_14;
  wire       [1:0]    CICC1851_mainAddrOne_15;
  wire       [11:0]   CICC1851_counterAddrTwo_15;
  wire       [11:0]   CICC1851_counterAddrTwo_16;
  wire       [11:0]   CICC1851_counterAddrTwo_17;
  wire       [1:0]    CICC1851_counterAddrTwo_18;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l664;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l664_1;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l664_2;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l665;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l665_1;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l665_2;
  reg                 inpDone;
  wire                when_SuperResolutionPart1_l79;
  reg                 startIn_regNext;
  wire                when_SuperResolutionPart1_l79_1;
  reg                 readDone;
  wire                when_SuperResolutionPart1_l82;
  reg                 startRead;
  wire                when_SuperResolutionPart1_l85;
  wire                when_SuperResolutionPart1_l85_1;
  reg                 slaveStart;
  wire                pixelsIn_fire;
  wire                when_SuperResolutionPart1_l88;
  wire                when_SuperResolutionPart1_l88_1;
  reg                 frameStart;
  reg        [7:0]    inpThreshold;
  reg        [9:0]    bmpWidth;
  reg        [9:0]    bmpHeight;
  reg                 holdBuffer;
  wire                when_SuperResolutionPart1_l103;
  reg                 writeDone;
  wire                when_SuperResolutionPart1_l106;
  reg                 bufferRowCount_willIncrement;
  reg                 bufferRowCount_willClear;
  reg        [9:0]    bufferRowCount_valueNext;
  reg        [9:0]    bufferRowCount_value;
  wire                bufferRowCount_willOverflowIfInc;
  wire                bufferRowCount_willOverflow;
  reg                 bufferEnable;
  wire                when_SuperResolutionPart1_l112;
  wire                when_SuperResolutionPart1_l112_1;
  reg                 bufferSwitch;
  wire                when_SuperResolutionPart1_l115;
  reg                 nextRowBuffer;
  wire                when_SuperResolutionPart1_l118;
  reg                 bufferReuse;
  reg                 bufferWAddr_willIncrement;
  reg                 bufferWAddr_willClear;
  reg        [9:0]    bufferWAddr_valueNext;
  reg        [9:0]    bufferWAddr_value;
  wire                bufferWAddr_willOverflowIfInc;
  wire                bufferWAddr_willOverflow;
  reg                 outPixelAddr_willIncrement;
  reg                 outPixelAddr_willClear;
  reg        [10:0]   outPixelAddr_valueNext;
  reg        [10:0]   outPixelAddr_value;
  wire                outPixelAddr_willOverflowIfInc;
  wire                outPixelAddr_willOverflow;
  reg                 outRowCount_willIncrement;
  reg                 outRowCount_willClear;
  reg        [10:0]   outRowCount_valueNext;
  reg        [10:0]   outRowCount_value;
  wire                outRowCount_willOverflowIfInc;
  wire                outRowCount_willOverflow;
  reg                 outReachRowEnd;
  reg                 outReachFinalRow;
  reg                 bufferReachRowEnd;
  reg                 bufferReachFinalRow;
  reg        [9:0]    mainAddrOne;
  reg        [9:0]    counterAddrOne;
  reg        [9:0]    mainAddrTwo;
  reg        [9:0]    counterAddrTwo;
  wire                validStream_valid;
  reg                 validStream_ready;
  wire                controlStream_valid;
  wire                controlStream_ready;
  wire                controlStream_payload_frameStart;
  wire                controlStream_payload_rowEnd;
  wire                controlStream_payload_passMode;
  wire                controlStream_payload_passValid;
  wire       [2:0]    controlStream_payload_onceMode;
  wire                controlStream_payload_onceValid;
  wire                controlStream_payload_mainCompare;
  wire                controlStream_payload_counterCompare;
  wire       [7:0]    controlStream_payload_mainDiff;
  wire       [7:0]    controlStream_payload_counterDiff;
  wire                controlStream_payload_twiceCompValid;
  wire       [2:0]    controlStream_payload_twiceMode;
  reg                 controls_frameStart;
  reg                 controls_rowEnd;
  reg                 controls_passMode;
  reg                 controls_passValid;
  reg        [2:0]    controls_onceMode;
  reg                 controls_onceValid;
  wire                controls_mainCompare;
  wire                controls_counterCompare;
  wire       [7:0]    controls_mainDiff;
  wire       [7:0]    controls_counterDiff;
  reg                 controls_twiceCompValid;
  reg        [2:0]    controls_twiceMode;
  wire       [29:0]   CICC1851_controls_frameStart;
  wire                mainAddrOneStream_valid;
  wire                mainAddrOneStream_ready;
  wire       [9:0]    mainAddrOneStream_payload;
  wire                counterAddrOneStream_valid;
  wire                counterAddrOneStream_ready;
  wire       [9:0]    counterAddrOneStream_payload;
  wire                mainAddrTwoStream_valid;
  wire                mainAddrTwoStream_ready;
  wire       [9:0]    mainAddrTwoStream_payload;
  wire                counterAddrTwoStream_valid;
  wire                counterAddrTwoStream_ready;
  wire       [9:0]    counterAddrTwoStream_payload;
  wire                mainAddrOneStream_s2mPipe_valid;
  reg                 mainAddrOneStream_s2mPipe_ready;
  wire       [9:0]    mainAddrOneStream_s2mPipe_payload;
  reg                 mainAddrOneStream_rValid;
  reg        [9:0]    mainAddrOneStream_rData;
  wire                mainAddrOneStream_s2mPipe_m2sPipe_valid;
  wire                mainAddrOneStream_s2mPipe_m2sPipe_ready;
  wire       [9:0]    mainAddrOneStream_s2mPipe_m2sPipe_payload;
  reg                 mainAddrOneStream_s2mPipe_rValid;
  reg        [9:0]    mainAddrOneStream_s2mPipe_rData;
  wire                when_Stream_l368;
  wire                CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_mainOnePixelStream_payload;
  reg                 CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_1;
  reg                 CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_mainOnePixelStream_payload_1;
  wire                readStage_mainOnePixelStream_valid;
  wire                readStage_mainOnePixelStream_ready;
  wire       [7:0]    readStage_mainOnePixelStream_payload;
  reg                 CICC1851_readStage_mainOnePixelStream_valid;
  reg        [7:0]    CICC1851_readStage_mainOnePixelStream_payload_2;
  wire                when_Stream_l368_1;
  wire                counterAddrOneStream_s2mPipe_valid;
  reg                 counterAddrOneStream_s2mPipe_ready;
  wire       [9:0]    counterAddrOneStream_s2mPipe_payload;
  reg                 counterAddrOneStream_rValid;
  reg        [9:0]    counterAddrOneStream_rData;
  wire                counterAddrOneStream_s2mPipe_m2sPipe_valid;
  wire                counterAddrOneStream_s2mPipe_m2sPipe_ready;
  wire       [9:0]    counterAddrOneStream_s2mPipe_m2sPipe_payload;
  reg                 counterAddrOneStream_s2mPipe_rValid;
  reg        [9:0]    counterAddrOneStream_s2mPipe_rData;
  wire                when_Stream_l368_2;
  wire                CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_counterOnePixelStream_payload;
  reg                 CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_2;
  reg                 CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_counterOnePixelStream_payload_1;
  wire                readStage_counterOnePixelStream_valid;
  wire                readStage_counterOnePixelStream_ready;
  wire       [7:0]    readStage_counterOnePixelStream_payload;
  reg                 CICC1851_readStage_counterOnePixelStream_valid;
  reg        [7:0]    CICC1851_readStage_counterOnePixelStream_payload_2;
  wire                when_Stream_l368_3;
  wire                mainAddrTwoStream_s2mPipe_valid;
  reg                 mainAddrTwoStream_s2mPipe_ready;
  wire       [9:0]    mainAddrTwoStream_s2mPipe_payload;
  reg                 mainAddrTwoStream_rValid;
  reg        [9:0]    mainAddrTwoStream_rData;
  wire                mainAddrTwoStream_s2mPipe_m2sPipe_valid;
  wire                mainAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire       [9:0]    mainAddrTwoStream_s2mPipe_m2sPipe_payload;
  reg                 mainAddrTwoStream_s2mPipe_rValid;
  reg        [9:0]    mainAddrTwoStream_s2mPipe_rData;
  wire                when_Stream_l368_4;
  wire                CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_mainTwoPixelStream_payload;
  reg                 CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_3;
  reg                 CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_mainTwoPixelStream_payload_1;
  wire                readStage_mainTwoPixelStream_valid;
  wire                readStage_mainTwoPixelStream_ready;
  wire       [7:0]    readStage_mainTwoPixelStream_payload;
  reg                 CICC1851_readStage_mainTwoPixelStream_valid;
  reg        [7:0]    CICC1851_readStage_mainTwoPixelStream_payload_2;
  wire                when_Stream_l368_5;
  wire                counterAddrTwoStream_s2mPipe_valid;
  reg                 counterAddrTwoStream_s2mPipe_ready;
  wire       [9:0]    counterAddrTwoStream_s2mPipe_payload;
  reg                 counterAddrTwoStream_rValid;
  reg        [9:0]    counterAddrTwoStream_rData;
  wire                counterAddrTwoStream_s2mPipe_m2sPipe_valid;
  wire                counterAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire       [9:0]    counterAddrTwoStream_s2mPipe_m2sPipe_payload;
  reg                 counterAddrTwoStream_s2mPipe_rValid;
  reg        [9:0]    counterAddrTwoStream_s2mPipe_rData;
  wire                when_Stream_l368_6;
  wire                CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_counterTwoPixelStream_payload;
  reg                 CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_4;
  reg                 CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_counterTwoPixelStream_payload_1;
  wire                readStage_counterTwoPixelStream_valid;
  wire                readStage_counterTwoPixelStream_ready;
  wire       [7:0]    readStage_counterTwoPixelStream_payload;
  reg                 CICC1851_readStage_counterTwoPixelStream_valid;
  reg        [7:0]    CICC1851_readStage_counterTwoPixelStream_payload_2;
  wire                when_Stream_l368_7;
  wire                controlStream_s2mPipe_valid;
  reg                 controlStream_s2mPipe_ready;
  wire                controlStream_s2mPipe_payload_frameStart;
  wire                controlStream_s2mPipe_payload_rowEnd;
  wire                controlStream_s2mPipe_payload_passMode;
  wire                controlStream_s2mPipe_payload_passValid;
  wire       [2:0]    controlStream_s2mPipe_payload_onceMode;
  wire                controlStream_s2mPipe_payload_onceValid;
  wire                controlStream_s2mPipe_payload_mainCompare;
  wire                controlStream_s2mPipe_payload_counterCompare;
  wire       [7:0]    controlStream_s2mPipe_payload_mainDiff;
  wire       [7:0]    controlStream_s2mPipe_payload_counterDiff;
  wire                controlStream_s2mPipe_payload_twiceCompValid;
  wire       [2:0]    controlStream_s2mPipe_payload_twiceMode;
  reg                 controlStream_rValid;
  reg                 controlStream_rData_frameStart;
  reg                 controlStream_rData_rowEnd;
  reg                 controlStream_rData_passMode;
  reg                 controlStream_rData_passValid;
  reg        [2:0]    controlStream_rData_onceMode;
  reg                 controlStream_rData_onceValid;
  reg                 controlStream_rData_mainCompare;
  reg                 controlStream_rData_counterCompare;
  reg        [7:0]    controlStream_rData_mainDiff;
  reg        [7:0]    controlStream_rData_counterDiff;
  reg                 controlStream_rData_twiceCompValid;
  reg        [2:0]    controlStream_rData_twiceMode;
  wire                controlStream_s2mPipe_m2sPipe_valid;
  reg                 controlStream_s2mPipe_m2sPipe_ready;
  wire                controlStream_s2mPipe_m2sPipe_payload_frameStart;
  wire                controlStream_s2mPipe_m2sPipe_payload_rowEnd;
  wire                controlStream_s2mPipe_m2sPipe_payload_passMode;
  wire                controlStream_s2mPipe_m2sPipe_payload_passValid;
  wire       [2:0]    controlStream_s2mPipe_m2sPipe_payload_onceMode;
  wire                controlStream_s2mPipe_m2sPipe_payload_onceValid;
  wire                controlStream_s2mPipe_m2sPipe_payload_mainCompare;
  wire                controlStream_s2mPipe_m2sPipe_payload_counterCompare;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_payload_mainDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_payload_counterDiff;
  wire                controlStream_s2mPipe_m2sPipe_payload_twiceCompValid;
  wire       [2:0]    controlStream_s2mPipe_m2sPipe_payload_twiceMode;
  reg                 controlStream_s2mPipe_rValid;
  reg                 controlStream_s2mPipe_rData_frameStart;
  reg                 controlStream_s2mPipe_rData_rowEnd;
  reg                 controlStream_s2mPipe_rData_passMode;
  reg                 controlStream_s2mPipe_rData_passValid;
  reg        [2:0]    controlStream_s2mPipe_rData_onceMode;
  reg                 controlStream_s2mPipe_rData_onceValid;
  reg                 controlStream_s2mPipe_rData_mainCompare;
  reg                 controlStream_s2mPipe_rData_counterCompare;
  reg        [7:0]    controlStream_s2mPipe_rData_mainDiff;
  reg        [7:0]    controlStream_s2mPipe_rData_counterDiff;
  reg                 controlStream_s2mPipe_rData_twiceCompValid;
  reg        [2:0]    controlStream_s2mPipe_rData_twiceMode;
  wire                when_Stream_l368_8;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_valid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_ready;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_frameStart;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_rowEnd;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passMode;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passValid;
  wire       [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceMode;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceValid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainCompare;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterCompare;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDiff;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceCompValid;
  wire       [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceMode;
  reg                 controlStream_s2mPipe_m2sPipe_rValid;
  reg                 controlStream_s2mPipe_m2sPipe_rData_frameStart;
  reg                 controlStream_s2mPipe_m2sPipe_rData_rowEnd;
  reg                 controlStream_s2mPipe_m2sPipe_rData_passMode;
  reg                 controlStream_s2mPipe_m2sPipe_rData_passValid;
  reg        [2:0]    controlStream_s2mPipe_m2sPipe_rData_onceMode;
  reg                 controlStream_s2mPipe_m2sPipe_rData_onceValid;
  reg                 controlStream_s2mPipe_m2sPipe_rData_mainCompare;
  reg                 controlStream_s2mPipe_m2sPipe_rData_counterCompare;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_rData_mainDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_rData_counterDiff;
  reg                 controlStream_s2mPipe_m2sPipe_rData_twiceCompValid;
  reg        [2:0]    controlStream_s2mPipe_m2sPipe_rData_twiceMode;
  wire                when_Stream_l368_9;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_valid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_frameStart;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_rowEnd;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_passMode;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_passValid;
  wire       [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_onceMode;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_onceValid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainCompare;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterCompare;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterDiff;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_twiceCompValid;
  wire       [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_twiceMode;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_frameStart;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_rowEnd;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_passMode;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_passValid;
  reg        [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_onceMode;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_onceValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainCompare;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterCompare;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterDiff;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_twiceCompValid;
  reg        [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_twiceMode;
  wire                readStage_controlPipe_valid;
  wire                readStage_controlPipe_ready;
  wire                readStage_controlPipe_payload_frameStart;
  wire                readStage_controlPipe_payload_rowEnd;
  wire                readStage_controlPipe_payload_passMode;
  wire                readStage_controlPipe_payload_passValid;
  wire       [2:0]    readStage_controlPipe_payload_onceMode;
  wire                readStage_controlPipe_payload_onceValid;
  wire                readStage_controlPipe_payload_mainCompare;
  wire                readStage_controlPipe_payload_counterCompare;
  wire       [7:0]    readStage_controlPipe_payload_mainDiff;
  wire       [7:0]    readStage_controlPipe_payload_counterDiff;
  wire                readStage_controlPipe_payload_twiceCompValid;
  wire       [2:0]    readStage_controlPipe_payload_twiceMode;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_frameStart;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_rowEnd;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_passMode;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_passValid;
  reg        [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_onceMode;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_onceValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainCompare;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterCompare;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterDiff;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_twiceCompValid;
  reg        [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_twiceMode;
  wire                when_Stream_l368_10;
  wire                readStage_mainOnePixelStream_s2mPipe_valid;
  reg                 readStage_mainOnePixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_mainOnePixelStream_s2mPipe_payload;
  reg                 readStage_mainOnePixelStream_rValid;
  reg        [7:0]    readStage_mainOnePixelStream_rData;
  wire                compareStage_mainOnePixelStream_valid;
  wire                compareStage_mainOnePixelStream_ready;
  wire       [7:0]    compareStage_mainOnePixelStream_payload;
  reg                 readStage_mainOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_mainOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_11;
  wire                readStage_counterOnePixelStream_s2mPipe_valid;
  reg                 readStage_counterOnePixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_counterOnePixelStream_s2mPipe_payload;
  reg                 readStage_counterOnePixelStream_rValid;
  reg        [7:0]    readStage_counterOnePixelStream_rData;
  wire                compareStage_counterOnePixelStream_valid;
  wire                compareStage_counterOnePixelStream_ready;
  wire       [7:0]    compareStage_counterOnePixelStream_payload;
  reg                 readStage_counterOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_counterOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_12;
  wire                readStage_mainTwoPixelStream_s2mPipe_valid;
  reg                 readStage_mainTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_mainTwoPixelStream_s2mPipe_payload;
  reg                 readStage_mainTwoPixelStream_rValid;
  reg        [7:0]    readStage_mainTwoPixelStream_rData;
  wire                compareStage_mainTwoPixelStream_valid;
  wire                compareStage_mainTwoPixelStream_ready;
  wire       [7:0]    compareStage_mainTwoPixelStream_payload;
  reg                 readStage_mainTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_mainTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_13;
  wire                readStage_counterTwoPixelStream_s2mPipe_valid;
  reg                 readStage_counterTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_counterTwoPixelStream_s2mPipe_payload;
  reg                 readStage_counterTwoPixelStream_rValid;
  reg        [7:0]    readStage_counterTwoPixelStream_rData;
  wire                compareStage_counterTwoPixelStream_valid;
  wire                compareStage_counterTwoPixelStream_ready;
  wire       [7:0]    compareStage_counterTwoPixelStream_payload;
  reg                 readStage_counterTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_counterTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_14;
  reg                 CICC1851_readStage_controlPipe_translated_payload_mainCompare;
  reg                 CICC1851_readStage_controlPipe_translated_payload_counterCompare;
  wire                when_SuperResolutionPart1_l205;
  wire                when_SuperResolutionPart1_l209;
  wire                when_SuperResolutionPart1_l213;
  wire                when_SuperResolutionPart1_l217;
  wire                when_SuperResolutionPart1_l228;
  wire                when_SuperResolutionPart1_l230;
  wire                when_SuperResolutionPart1_l234;
  wire                when_SuperResolutionPart1_l236;
  wire                when_SuperResolutionPart1_l241;
  wire                when_SuperResolutionPart1_l246;
  wire                readStage_controlPipe_translated_valid;
  wire                readStage_controlPipe_translated_ready;
  wire                readStage_controlPipe_translated_payload_frameStart;
  wire                readStage_controlPipe_translated_payload_rowEnd;
  wire                readStage_controlPipe_translated_payload_passMode;
  wire                readStage_controlPipe_translated_payload_passValid;
  wire       [2:0]    readStage_controlPipe_translated_payload_onceMode;
  wire                readStage_controlPipe_translated_payload_onceValid;
  wire                readStage_controlPipe_translated_payload_mainCompare;
  wire                readStage_controlPipe_translated_payload_counterCompare;
  wire       [7:0]    readStage_controlPipe_translated_payload_mainDiff;
  wire       [7:0]    readStage_controlPipe_translated_payload_counterDiff;
  wire                readStage_controlPipe_translated_payload_twiceCompValid;
  wire       [2:0]    readStage_controlPipe_translated_payload_twiceMode;
  wire                readStage_controlPipe_translated_s2mPipe_valid;
  reg                 readStage_controlPipe_translated_s2mPipe_ready;
  wire                readStage_controlPipe_translated_s2mPipe_payload_frameStart;
  wire                readStage_controlPipe_translated_s2mPipe_payload_rowEnd;
  wire                readStage_controlPipe_translated_s2mPipe_payload_passMode;
  wire                readStage_controlPipe_translated_s2mPipe_payload_passValid;
  wire       [2:0]    readStage_controlPipe_translated_s2mPipe_payload_onceMode;
  wire                readStage_controlPipe_translated_s2mPipe_payload_onceValid;
  wire                readStage_controlPipe_translated_s2mPipe_payload_mainCompare;
  wire                readStage_controlPipe_translated_s2mPipe_payload_counterCompare;
  wire       [7:0]    readStage_controlPipe_translated_s2mPipe_payload_mainDiff;
  wire       [7:0]    readStage_controlPipe_translated_s2mPipe_payload_counterDiff;
  wire                readStage_controlPipe_translated_s2mPipe_payload_twiceCompValid;
  wire       [2:0]    readStage_controlPipe_translated_s2mPipe_payload_twiceMode;
  reg                 readStage_controlPipe_translated_rValid;
  reg                 readStage_controlPipe_translated_rData_frameStart;
  reg                 readStage_controlPipe_translated_rData_rowEnd;
  reg                 readStage_controlPipe_translated_rData_passMode;
  reg                 readStage_controlPipe_translated_rData_passValid;
  reg        [2:0]    readStage_controlPipe_translated_rData_onceMode;
  reg                 readStage_controlPipe_translated_rData_onceValid;
  reg                 readStage_controlPipe_translated_rData_mainCompare;
  reg                 readStage_controlPipe_translated_rData_counterCompare;
  reg        [7:0]    readStage_controlPipe_translated_rData_mainDiff;
  reg        [7:0]    readStage_controlPipe_translated_rData_counterDiff;
  reg                 readStage_controlPipe_translated_rData_twiceCompValid;
  reg        [2:0]    readStage_controlPipe_translated_rData_twiceMode;
  wire                compareStage_controlPipe_valid;
  wire                compareStage_controlPipe_ready;
  wire                compareStage_controlPipe_payload_frameStart;
  wire                compareStage_controlPipe_payload_rowEnd;
  wire                compareStage_controlPipe_payload_passMode;
  wire                compareStage_controlPipe_payload_passValid;
  wire       [2:0]    compareStage_controlPipe_payload_onceMode;
  wire                compareStage_controlPipe_payload_onceValid;
  wire                compareStage_controlPipe_payload_mainCompare;
  wire                compareStage_controlPipe_payload_counterCompare;
  wire       [7:0]    compareStage_controlPipe_payload_mainDiff;
  wire       [7:0]    compareStage_controlPipe_payload_counterDiff;
  wire                compareStage_controlPipe_payload_twiceCompValid;
  wire       [2:0]    compareStage_controlPipe_payload_twiceMode;
  reg                 readStage_controlPipe_translated_s2mPipe_rValid;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_frameStart;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_rowEnd;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_passMode;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_passValid;
  reg        [2:0]    readStage_controlPipe_translated_s2mPipe_rData_onceMode;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_onceValid;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_mainCompare;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_counterCompare;
  reg        [7:0]    readStage_controlPipe_translated_s2mPipe_rData_mainDiff;
  reg        [7:0]    readStage_controlPipe_translated_s2mPipe_rData_counterDiff;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_twiceCompValid;
  reg        [2:0]    readStage_controlPipe_translated_s2mPipe_rData_twiceMode;
  wire                when_Stream_l368_15;
  wire                compareStage_mainOnePixelStream_s2mPipe_valid;
  reg                 compareStage_mainOnePixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_mainOnePixelStream_s2mPipe_payload;
  reg                 compareStage_mainOnePixelStream_rValid;
  reg        [7:0]    compareStage_mainOnePixelStream_rData;
  wire                diffStage_mainOnePixelStream_valid;
  wire                diffStage_mainOnePixelStream_ready;
  wire       [7:0]    diffStage_mainOnePixelStream_payload;
  reg                 compareStage_mainOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_mainOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_16;
  wire                compareStage_counterOnePixelStream_s2mPipe_valid;
  reg                 compareStage_counterOnePixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_counterOnePixelStream_s2mPipe_payload;
  reg                 compareStage_counterOnePixelStream_rValid;
  reg        [7:0]    compareStage_counterOnePixelStream_rData;
  wire                diffStage_counterOnePixelStream_valid;
  wire                diffStage_counterOnePixelStream_ready;
  wire       [7:0]    diffStage_counterOnePixelStream_payload;
  reg                 compareStage_counterOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_counterOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_17;
  wire                compareStage_mainTwoPixelStream_s2mPipe_valid;
  reg                 compareStage_mainTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_mainTwoPixelStream_s2mPipe_payload;
  reg                 compareStage_mainTwoPixelStream_rValid;
  reg        [7:0]    compareStage_mainTwoPixelStream_rData;
  wire                diffStage_mainTwoPixelStream_valid;
  wire                diffStage_mainTwoPixelStream_ready;
  wire       [7:0]    diffStage_mainTwoPixelStream_payload;
  reg                 compareStage_mainTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_mainTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_18;
  wire                compareStage_counterTwoPixelStream_s2mPipe_valid;
  reg                 compareStage_counterTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_counterTwoPixelStream_s2mPipe_payload;
  reg                 compareStage_counterTwoPixelStream_rValid;
  reg        [7:0]    compareStage_counterTwoPixelStream_rData;
  wire                diffStage_counterTwoPixelStream_valid;
  wire                diffStage_counterTwoPixelStream_ready;
  wire       [7:0]    diffStage_counterTwoPixelStream_payload;
  reg                 compareStage_counterTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_counterTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_19;
  reg        [7:0]    CICC1851_compareStage_controlPipe_translated_payload_mainDiff;
  reg        [7:0]    CICC1851_compareStage_controlPipe_translated_payload_counterDiff;
  wire                compareStage_controlPipe_translated_valid;
  wire                compareStage_controlPipe_translated_ready;
  wire                compareStage_controlPipe_translated_payload_frameStart;
  wire                compareStage_controlPipe_translated_payload_rowEnd;
  wire                compareStage_controlPipe_translated_payload_passMode;
  wire                compareStage_controlPipe_translated_payload_passValid;
  wire       [2:0]    compareStage_controlPipe_translated_payload_onceMode;
  wire                compareStage_controlPipe_translated_payload_onceValid;
  wire                compareStage_controlPipe_translated_payload_mainCompare;
  wire                compareStage_controlPipe_translated_payload_counterCompare;
  wire       [7:0]    compareStage_controlPipe_translated_payload_mainDiff;
  wire       [7:0]    compareStage_controlPipe_translated_payload_counterDiff;
  wire                compareStage_controlPipe_translated_payload_twiceCompValid;
  wire       [2:0]    compareStage_controlPipe_translated_payload_twiceMode;
  wire                compareStage_controlPipe_translated_s2mPipe_valid;
  reg                 compareStage_controlPipe_translated_s2mPipe_ready;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_frameStart;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_rowEnd;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_passMode;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_passValid;
  wire       [2:0]    compareStage_controlPipe_translated_s2mPipe_payload_onceMode;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_onceValid;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_mainCompare;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_counterCompare;
  wire       [7:0]    compareStage_controlPipe_translated_s2mPipe_payload_mainDiff;
  wire       [7:0]    compareStage_controlPipe_translated_s2mPipe_payload_counterDiff;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_twiceCompValid;
  wire       [2:0]    compareStage_controlPipe_translated_s2mPipe_payload_twiceMode;
  reg                 compareStage_controlPipe_translated_rValid;
  reg                 compareStage_controlPipe_translated_rData_frameStart;
  reg                 compareStage_controlPipe_translated_rData_rowEnd;
  reg                 compareStage_controlPipe_translated_rData_passMode;
  reg                 compareStage_controlPipe_translated_rData_passValid;
  reg        [2:0]    compareStage_controlPipe_translated_rData_onceMode;
  reg                 compareStage_controlPipe_translated_rData_onceValid;
  reg                 compareStage_controlPipe_translated_rData_mainCompare;
  reg                 compareStage_controlPipe_translated_rData_counterCompare;
  reg        [7:0]    compareStage_controlPipe_translated_rData_mainDiff;
  reg        [7:0]    compareStage_controlPipe_translated_rData_counterDiff;
  reg                 compareStage_controlPipe_translated_rData_twiceCompValid;
  reg        [2:0]    compareStage_controlPipe_translated_rData_twiceMode;
  wire                diffStage_controlPipe_valid;
  wire                diffStage_controlPipe_ready;
  wire                diffStage_controlPipe_payload_frameStart;
  wire                diffStage_controlPipe_payload_rowEnd;
  wire                diffStage_controlPipe_payload_passMode;
  wire                diffStage_controlPipe_payload_passValid;
  wire       [2:0]    diffStage_controlPipe_payload_onceMode;
  wire                diffStage_controlPipe_payload_onceValid;
  wire                diffStage_controlPipe_payload_mainCompare;
  wire                diffStage_controlPipe_payload_counterCompare;
  wire       [7:0]    diffStage_controlPipe_payload_mainDiff;
  wire       [7:0]    diffStage_controlPipe_payload_counterDiff;
  wire                diffStage_controlPipe_payload_twiceCompValid;
  wire       [2:0]    diffStage_controlPipe_payload_twiceMode;
  reg                 compareStage_controlPipe_translated_s2mPipe_rValid;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_frameStart;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_rowEnd;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_passMode;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_passValid;
  reg        [2:0]    compareStage_controlPipe_translated_s2mPipe_rData_onceMode;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_onceValid;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_mainCompare;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_counterCompare;
  reg        [7:0]    compareStage_controlPipe_translated_s2mPipe_rData_mainDiff;
  reg        [7:0]    compareStage_controlPipe_translated_s2mPipe_rData_counterDiff;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_twiceCompValid;
  reg        [2:0]    compareStage_controlPipe_translated_s2mPipe_rData_twiceMode;
  wire                when_Stream_l368_20;
  wire                diffStage_mainOnePixelStream_s2mPipe_valid;
  reg                 diffStage_mainOnePixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_mainOnePixelStream_s2mPipe_payload;
  reg                 diffStage_mainOnePixelStream_rValid;
  reg        [7:0]    diffStage_mainOnePixelStream_rData;
  wire                resultStage_mainOnePixelStream_valid;
  wire                resultStage_mainOnePixelStream_ready;
  wire       [7:0]    resultStage_mainOnePixelStream_payload;
  reg                 diffStage_mainOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_mainOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_21;
  wire                diffStage_counterOnePixelStream_s2mPipe_valid;
  reg                 diffStage_counterOnePixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_counterOnePixelStream_s2mPipe_payload;
  reg                 diffStage_counterOnePixelStream_rValid;
  reg        [7:0]    diffStage_counterOnePixelStream_rData;
  wire                resultStage_counterOnePixelStream_valid;
  wire                resultStage_counterOnePixelStream_ready;
  wire       [7:0]    resultStage_counterOnePixelStream_payload;
  reg                 diffStage_counterOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_counterOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_22;
  wire                diffStage_mainTwoPixelStream_s2mPipe_valid;
  reg                 diffStage_mainTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_mainTwoPixelStream_s2mPipe_payload;
  reg                 diffStage_mainTwoPixelStream_rValid;
  reg        [7:0]    diffStage_mainTwoPixelStream_rData;
  wire                resultStage_mainTwoPixelStream_valid;
  wire                resultStage_mainTwoPixelStream_ready;
  wire       [7:0]    resultStage_mainTwoPixelStream_payload;
  reg                 diffStage_mainTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_mainTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_23;
  wire                diffStage_counterTwoPixelStream_s2mPipe_valid;
  reg                 diffStage_counterTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_counterTwoPixelStream_s2mPipe_payload;
  reg                 diffStage_counterTwoPixelStream_rValid;
  reg        [7:0]    diffStage_counterTwoPixelStream_rData;
  wire                resultStage_counterTwoPixelStream_valid;
  wire                resultStage_counterTwoPixelStream_ready;
  wire       [7:0]    resultStage_counterTwoPixelStream_payload;
  reg                 diffStage_counterTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_counterTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_24;
  wire                diffStage_controlPipe_fork_io_outputs_0_s2mPipe_valid;
  reg                 diffStage_controlPipe_fork_io_outputs_0_s2mPipe_ready;
  wire                diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_frameStart;
  wire                diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_rowEnd;
  wire                diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_passMode;
  wire                diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_passValid;
  wire       [2:0]    diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_onceMode;
  wire                diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_onceValid;
  wire                diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_mainCompare;
  wire                diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_counterCompare;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_mainDiff;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_counterDiff;
  wire                diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_twiceCompValid;
  wire       [2:0]    diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_twiceMode;
  reg                 diffStage_controlPipe_fork_io_outputs_0_rValid;
  reg                 diffStage_controlPipe_fork_io_outputs_0_rData_frameStart;
  reg                 diffStage_controlPipe_fork_io_outputs_0_rData_rowEnd;
  reg                 diffStage_controlPipe_fork_io_outputs_0_rData_passMode;
  reg                 diffStage_controlPipe_fork_io_outputs_0_rData_passValid;
  reg        [2:0]    diffStage_controlPipe_fork_io_outputs_0_rData_onceMode;
  reg                 diffStage_controlPipe_fork_io_outputs_0_rData_onceValid;
  reg                 diffStage_controlPipe_fork_io_outputs_0_rData_mainCompare;
  reg                 diffStage_controlPipe_fork_io_outputs_0_rData_counterCompare;
  reg        [7:0]    diffStage_controlPipe_fork_io_outputs_0_rData_mainDiff;
  reg        [7:0]    diffStage_controlPipe_fork_io_outputs_0_rData_counterDiff;
  reg                 diffStage_controlPipe_fork_io_outputs_0_rData_twiceCompValid;
  reg        [2:0]    diffStage_controlPipe_fork_io_outputs_0_rData_twiceMode;
  wire                resultStage_controlPipe_valid;
  wire                resultStage_controlPipe_ready;
  wire                resultStage_controlPipe_payload_frameStart;
  wire                resultStage_controlPipe_payload_rowEnd;
  wire                resultStage_controlPipe_payload_passMode;
  wire                resultStage_controlPipe_payload_passValid;
  wire       [2:0]    resultStage_controlPipe_payload_onceMode;
  wire                resultStage_controlPipe_payload_onceValid;
  wire                resultStage_controlPipe_payload_mainCompare;
  wire                resultStage_controlPipe_payload_counterCompare;
  wire       [7:0]    resultStage_controlPipe_payload_mainDiff;
  wire       [7:0]    resultStage_controlPipe_payload_counterDiff;
  wire                resultStage_controlPipe_payload_twiceCompValid;
  wire       [2:0]    resultStage_controlPipe_payload_twiceMode;
  reg                 diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rValid;
  reg                 diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_frameStart;
  reg                 diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_rowEnd;
  reg                 diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_passMode;
  reg                 diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_passValid;
  reg        [2:0]    diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_onceMode;
  reg                 diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_onceValid;
  reg                 diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_mainCompare;
  reg                 diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_counterCompare;
  reg        [7:0]    diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_mainDiff;
  reg        [7:0]    diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_counterDiff;
  reg                 diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_twiceCompValid;
  reg        [2:0]    diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_twiceMode;
  wire                when_Stream_l368_25;
  wire                resultStage_pixelStream_valid;
  wire                resultStage_pixelStream_ready;
  reg        [7:0]    resultStage_pixelStream_payload;
  wire                when_SuperResolutionPart1_l339;
  wire                when_SuperResolutionPart1_l343;
  wire                when_SuperResolutionPart1_l347;
  wire                when_SuperResolutionPart1_l351;
  wire                when_SuperResolutionPart1_l362;
  wire                when_SuperResolutionPart1_l363;
  wire                when_SuperResolutionPart1_l366;
  wire                when_SuperResolutionPart1_l371;
  wire                when_SuperResolutionPart1_l372;
  wire                when_SuperResolutionPart1_l375;
  wire                when_SuperResolutionPart1_l381;
  wire                when_SuperResolutionPart1_l386;
  wire                resultStage_pixelStream_s2mPipe_valid;
  reg                 resultStage_pixelStream_s2mPipe_ready;
  wire       [7:0]    resultStage_pixelStream_s2mPipe_payload;
  reg                 resultStage_pixelStream_rValid;
  reg        [7:0]    resultStage_pixelStream_rData;
  wire                resultStage_resultStream_valid;
  wire                resultStage_resultStream_ready;
  wire       [7:0]    resultStage_resultStream_payload;
  reg                 resultStage_pixelStream_s2mPipe_rValid;
  reg        [7:0]    resultStage_pixelStream_s2mPipe_rData;
  wire                when_Stream_l368_26;
  wire                CICC1851_resultStage_mainOnePixelStream_ready;
  reg                 CICC1851_resultStage_mainOnePixelStream_ready_1;
  wire                CICC1851_resultStage_mainOnePixelStream_ready_2;
  wire                when_Stream_l438;
  reg                 resultsJoin_valid;
  wire                resultsJoin_ready;
  wire                pixelsStream_valid;
  wire                pixelsStream_ready;
  wire       [7:0]    pixelsStream_payload_pixel;
  wire                pixelsStream_payload_frameStart;
  wire                pixelsStream_payload_rowEnd;
  wire                pixelsStream_s2mPipe_valid;
  reg                 pixelsStream_s2mPipe_ready;
  wire       [7:0]    pixelsStream_s2mPipe_payload_pixel;
  wire                pixelsStream_s2mPipe_payload_frameStart;
  wire                pixelsStream_s2mPipe_payload_rowEnd;
  reg                 pixelsStream_rValid;
  reg        [7:0]    pixelsStream_rData_pixel;
  reg                 pixelsStream_rData_frameStart;
  reg                 pixelsStream_rData_rowEnd;
  wire                pixelsStream_s2mPipe_m2sPipe_valid;
  wire                pixelsStream_s2mPipe_m2sPipe_ready;
  wire       [7:0]    pixelsStream_s2mPipe_m2sPipe_payload_pixel;
  wire                pixelsStream_s2mPipe_m2sPipe_payload_frameStart;
  wire                pixelsStream_s2mPipe_m2sPipe_payload_rowEnd;
  reg                 pixelsStream_s2mPipe_rValid;
  reg        [7:0]    pixelsStream_s2mPipe_rData_pixel;
  reg                 pixelsStream_s2mPipe_rData_frameStart;
  reg                 pixelsStream_s2mPipe_rData_rowEnd;
  wire                when_Stream_l368_27;
  wire                pixelsIn_s2mPipe_valid;
  reg                 pixelsIn_s2mPipe_ready;
  wire       [7:0]    pixelsIn_s2mPipe_payload_pixel;
  wire                pixelsIn_s2mPipe_payload_frameStart;
  wire                pixelsIn_s2mPipe_payload_rowEnd;
  reg                 pixelsIn_rValid;
  reg        [7:0]    pixelsIn_rData_pixel;
  reg                 pixelsIn_rData_frameStart;
  reg                 pixelsIn_rData_rowEnd;
  wire                pixelsIn_s2mPipe_m2sPipe_valid;
  wire                pixelsIn_s2mPipe_m2sPipe_ready;
  wire       [7:0]    pixelsIn_s2mPipe_m2sPipe_payload_pixel;
  wire                pixelsIn_s2mPipe_m2sPipe_payload_frameStart;
  wire                pixelsIn_s2mPipe_m2sPipe_payload_rowEnd;
  reg                 pixelsIn_s2mPipe_rValid;
  reg        [7:0]    pixelsIn_s2mPipe_rData_pixel;
  reg                 pixelsIn_s2mPipe_rData_frameStart;
  reg                 pixelsIn_s2mPipe_rData_rowEnd;
  wire                when_Stream_l368_28;
  wire                passPixels_valid;
  wire                passPixels_ready;
  wire       [7:0]    passPixels_payload_pixel;
  wire                passPixels_payload_frameStart;
  wire                passPixels_payload_rowEnd;
  wire                passPixels_fire;
  wire                when_SuperResolutionPart1_l421;
  wire                passPixels_fire_1;
  wire                when_SuperResolutionPart1_l422;
  wire                passPixels_fire_2;
  wire                when_SuperResolutionPart1_l425;
  wire                passPixels_fire_3;
  wire                when_SuperResolutionPart1_l438;
  wire                passPixels_fire_4;
  wire                when_SuperResolutionPart1_l439;
  wire                when_SuperResolutionPart1_l442;
  wire                controlStream_fire;
  wire                when_SuperResolutionPart1_l447;
  wire                when_SuperResolutionPart1_l449;
  wire                passPixels_fire_5;
  wire                when_SuperResolutionPart1_l453;
  wire                passPixels_fire_6;
  wire                passPixels_fire_7;
  wire                passPixels_fire_8;
  wire                controlStateMachine_wantExit;
  reg                 controlStateMachine_wantStart;
  wire                controlStateMachine_wantKill;
  reg        [2:0]    controlStateMachine_stateReg;
  reg        [2:0]    controlStateMachine_stateNext;
  wire                when_SuperResolutionPart1_l482;
  wire                passPixels_fire_9;
  wire                when_SuperResolutionPart1_l484;
  wire                passPixels_fire_10;
  wire                when_SuperResolutionPart1_l489;
  wire                controlStream_fire_1;
  wire                when_SuperResolutionPart1_l498;
  wire                passPixels_fire_11;
  wire                when_SuperResolutionPart1_l500;
  wire                controlStream_fire_2;
  wire                when_SuperResolutionPart1_l507;
  wire                controlStream_fire_3;
  wire                when_SuperResolutionPart1_l510;
  wire                controlStream_fire_4;
  wire                when_SuperResolutionPart1_l511;
  wire                controlStream_fire_5;
  wire                when_SuperResolutionPart1_l513;
  wire                controlStream_fire_6;
  wire                when_SuperResolutionPart1_l537;
  wire                controlStream_fire_7;
  wire                when_SuperResolutionPart1_l542;
  wire                controlStream_fire_8;
  wire                passPixels_fire_12;
  wire                when_SuperResolutionPart1_l563;
  wire                controlStream_fire_9;
  wire                when_SuperResolutionPart1_l578;
  wire                controlStream_fire_10;
  wire                when_SuperResolutionPart1_l579;
  wire                controlStream_fire_11;
  wire                when_SuperResolutionPart1_l581;
  wire                controlStream_fire_12;
  wire                controlStream_fire_13;
  wire                when_SuperResolutionPart1_l612;
  wire                controlStream_fire_14;
  wire                when_SuperResolutionPart1_l664;
  wire                controlStream_fire_15;
  wire                when_SuperResolutionPart1_l665;
  wire                controlStream_fire_16;
  wire                when_SuperResolutionPart1_l667;
  wire                controlStream_fire_17;
  `ifndef SYNTHESIS
  reg [39:0] controlStateMachine_stateReg_string;
  reg [39:0] controlStateMachine_stateNext_string;
  `endif

  reg [7:0] lineBufferOne [0:959];
  reg [7:0] lineBufferTwo [0:959];

  assign CICC1851_bufferRowCount_valueNext_1 = bufferRowCount_willIncrement;
  assign CICC1851_bufferRowCount_valueNext = {9'd0, CICC1851_bufferRowCount_valueNext_1};
  assign CICC1851_bufferWAddr_valueNext_1 = bufferWAddr_willIncrement;
  assign CICC1851_bufferWAddr_valueNext = {9'd0, CICC1851_bufferWAddr_valueNext_1};
  assign CICC1851_outPixelAddr_valueNext_1 = outPixelAddr_willIncrement;
  assign CICC1851_outPixelAddr_valueNext = {10'd0, CICC1851_outPixelAddr_valueNext_1};
  assign CICC1851_outRowCount_valueNext_1 = outRowCount_willIncrement;
  assign CICC1851_outRowCount_valueNext = {10'd0, CICC1851_outRowCount_valueNext_1};
  assign CICC1851_mainAddrOne = (outPixelAddr_value / 2'b10);
  assign CICC1851_counterAddrOne = (outPixelAddr_value / 2'b10);
  assign CICC1851_mainAddrTwo = (outPixelAddr_value / 2'b10);
  assign CICC1851_counterAddrTwo = (outPixelAddr_value / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload = (CICC1851_resultStage_pixelStream_payload_1 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_1 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_2 = (CICC1851_resultStage_pixelStream_payload_3 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_3 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_4 = (CICC1851_resultStage_pixelStream_payload_5 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_5 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_mainTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_6 = (CICC1851_resultStage_pixelStream_payload_7 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_7 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_mainOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_8 = (CICC1851_resultStage_pixelStream_payload_9 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_9 = ({1'b0,diffStage_counterOnePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_10 = (CICC1851_resultStage_pixelStream_payload_11 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_11 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_mainTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_12 = (CICC1851_resultStage_pixelStream_payload_13 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_13 = ({1'b0,diffStage_counterOnePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_14 = (CICC1851_resultStage_pixelStream_payload_15 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_15 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_mainTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_16 = (CICC1851_resultStage_pixelStream_payload_17 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_17 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_18 = (CICC1851_resultStage_pixelStream_payload_19 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_19 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_when_SuperResolutionPart1_l421 = (bmpWidth - 10'h002);
  assign CICC1851_when_SuperResolutionPart1_l422 = (bmpHeight - 10'h002);
  assign CICC1851_when_SuperResolutionPart1_l447 = (outRowCount_value % 2'b10);
  assign CICC1851_when_SuperResolutionPart1_l482 = (outRowCount_value % 2'b10);
  assign CICC1851_when_SuperResolutionPart1_l484 = (outPixelAddr_value % 2'b10);
  assign CICC1851_when_SuperResolutionPart1_l489 = (outPixelAddr_value % 2'b10);
  assign CICC1851_when_SuperResolutionPart1_l498 = {1'd0, outRowCount_value};
  assign CICC1851_when_SuperResolutionPart1_l498_1 = (2'b10 * bufferRowCount_value);
  assign CICC1851_when_SuperResolutionPart1_l500 = (2'b10 * bufferWAddr_value);
  assign CICC1851_when_SuperResolutionPart1_l500_1 = ({1'b0,outPixelAddr_value} + CICC1851_when_SuperResolutionPart1_l500_2);
  assign CICC1851_when_SuperResolutionPart1_l500_3 = {1'b0,2'b10};
  assign CICC1851_when_SuperResolutionPart1_l500_2 = {9'd0, CICC1851_when_SuperResolutionPart1_l500_3};
  assign CICC1851_when_SuperResolutionPart1_l510 = {1'd0, outPixelAddr_value};
  assign CICC1851_when_SuperResolutionPart1_l510_1 = (CICC1851_when_SuperResolutionPart1_l510_2 - 12'h002);
  assign CICC1851_when_SuperResolutionPart1_l510_2 = (2'b10 * bmpWidth);
  assign CICC1851_when_SuperResolutionPart1_l511 = {1'd0, outRowCount_value};
  assign CICC1851_when_SuperResolutionPart1_l511_1 = (CICC1851_when_SuperResolutionPart1_l511_2 - 12'h002);
  assign CICC1851_when_SuperResolutionPart1_l511_2 = (2'b10 * bmpHeight);
  assign CICC1851_when_SuperResolutionPart1_l537 = (outRowCount_value % 2'b10);
  assign CICC1851_when_SuperResolutionPart1_l542_1 = (11'h002 + outRowCount_value);
  assign CICC1851_when_SuperResolutionPart1_l542 = {1'd0, CICC1851_when_SuperResolutionPart1_l542_1};
  assign CICC1851_when_SuperResolutionPart1_l542_2 = (2'b10 * bufferRowCount_value);
  assign CICC1851_mainAddrOne_1 = (CICC1851_mainAddrOne_2 / 2'b10);
  assign CICC1851_mainAddrOne_2 = (outPixelAddr_value - 11'h001);
  assign CICC1851_counterAddrOne_1 = (CICC1851_counterAddrOne_2 / 2'b10);
  assign CICC1851_counterAddrOne_2 = (outPixelAddr_value - 11'h001);
  assign CICC1851_counterAddrOne_3 = (CICC1851_counterAddrOne_4 / 2'b10);
  assign CICC1851_counterAddrOne_4 = ({1'b0,outPixelAddr_value} + CICC1851_counterAddrOne_5);
  assign CICC1851_counterAddrOne_6 = {1'b0,1'b1};
  assign CICC1851_counterAddrOne_5 = {10'd0, CICC1851_counterAddrOne_6};
  assign CICC1851_controls_onceMode = 1'b1;
  assign CICC1851_mainAddrTwo_1 = (CICC1851_mainAddrTwo_2 / 2'b10);
  assign CICC1851_mainAddrTwo_2 = (outPixelAddr_value - 11'h001);
  assign CICC1851_counterAddrTwo_1 = (CICC1851_counterAddrTwo_2 / 2'b10);
  assign CICC1851_counterAddrTwo_2 = (outPixelAddr_value - 11'h001);
  assign CICC1851_counterAddrTwo_3 = (CICC1851_counterAddrTwo_4 / 2'b10);
  assign CICC1851_counterAddrTwo_4 = ({1'b0,outPixelAddr_value} + CICC1851_counterAddrTwo_5);
  assign CICC1851_counterAddrTwo_6 = {1'b0,1'b1};
  assign CICC1851_counterAddrTwo_5 = {10'd0, CICC1851_counterAddrTwo_6};
  assign CICC1851_when_SuperResolutionPart1_l563 = (2'b10 * bufferWAddr_value);
  assign CICC1851_when_SuperResolutionPart1_l563_1 = ({1'b0,outPixelAddr_value} + CICC1851_when_SuperResolutionPart1_l563_2);
  assign CICC1851_when_SuperResolutionPart1_l563_3 = {1'b0,2'b10};
  assign CICC1851_when_SuperResolutionPart1_l563_2 = {9'd0, CICC1851_when_SuperResolutionPart1_l563_3};
  assign CICC1851_controls_onceMode_1 = 2'b10;
  assign CICC1851_controls_onceMode_2 = 2'b11;
  assign CICC1851_mainAddrOne_3 = (outPixelAddr_value / 2'b10);
  assign CICC1851_mainAddrTwo_3 = (outPixelAddr_value / 2'b10);
  assign CICC1851_when_SuperResolutionPart1_l578 = {1'd0, outPixelAddr_value};
  assign CICC1851_when_SuperResolutionPart1_l578_1 = (CICC1851_when_SuperResolutionPart1_l578_2 - 12'h002);
  assign CICC1851_when_SuperResolutionPart1_l578_2 = (2'b10 * bmpWidth);
  assign CICC1851_when_SuperResolutionPart1_l579 = {1'd0, outRowCount_value};
  assign CICC1851_when_SuperResolutionPart1_l579_1 = (CICC1851_when_SuperResolutionPart1_l579_2 - 12'h002);
  assign CICC1851_when_SuperResolutionPart1_l579_2 = (2'b10 * bmpHeight);
  assign CICC1851_mainAddrOne_4 = (CICC1851_mainAddrOne_5 / 2'b10);
  assign CICC1851_mainAddrOne_5 = (outPixelAddr_value - 11'h001);
  assign CICC1851_mainAddrOne_6 = (CICC1851_mainAddrOne_7 / 2'b10);
  assign CICC1851_mainAddrOne_7 = (outPixelAddr_value - 11'h001);
  assign CICC1851_counterAddrOne_7 = (CICC1851_counterAddrOne_8 / 2'b10);
  assign CICC1851_counterAddrOne_8 = ({1'b0,outPixelAddr_value} + CICC1851_counterAddrOne_9);
  assign CICC1851_counterAddrOne_10 = {1'b0,1'b1};
  assign CICC1851_counterAddrOne_9 = {10'd0, CICC1851_counterAddrOne_10};
  assign CICC1851_mainAddrTwo_4 = (CICC1851_mainAddrTwo_5 / 2'b10);
  assign CICC1851_mainAddrTwo_5 = (outPixelAddr_value - 11'h001);
  assign CICC1851_mainAddrTwo_6 = (CICC1851_mainAddrTwo_7 / 2'b10);
  assign CICC1851_mainAddrTwo_7 = (outPixelAddr_value - 11'h001);
  assign CICC1851_counterAddrTwo_7 = (CICC1851_counterAddrTwo_8 / 2'b10);
  assign CICC1851_counterAddrTwo_8 = ({1'b0,outPixelAddr_value} + CICC1851_counterAddrTwo_9);
  assign CICC1851_counterAddrTwo_10 = {1'b0,1'b1};
  assign CICC1851_counterAddrTwo_9 = {10'd0, CICC1851_counterAddrTwo_10};
  assign CICC1851_mainAddrOne_8 = (CICC1851_mainAddrOne_9 / 2'b10);
  assign CICC1851_mainAddrOne_9 = (outPixelAddr_value - 11'h001);
  assign CICC1851_counterAddrTwo_11 = (CICC1851_counterAddrTwo_12 / 2'b10);
  assign CICC1851_counterAddrTwo_12 = (outPixelAddr_value - 11'h001);
  assign CICC1851_mainAddrTwo_8 = (CICC1851_mainAddrTwo_9 / 2'b10);
  assign CICC1851_mainAddrTwo_9 = (outPixelAddr_value - 11'h001);
  assign CICC1851_counterAddrOne_11 = (CICC1851_counterAddrOne_12 / 2'b10);
  assign CICC1851_counterAddrOne_12 = (outPixelAddr_value - 11'h001);
  assign CICC1851_mainAddrTwo_10 = (CICC1851_mainAddrTwo_11 / 2'b10);
  assign CICC1851_mainAddrTwo_11 = ({1'b0,outPixelAddr_value} + CICC1851_mainAddrTwo_12);
  assign CICC1851_mainAddrTwo_13 = {1'b0,1'b1};
  assign CICC1851_mainAddrTwo_12 = {10'd0, CICC1851_mainAddrTwo_13};
  assign CICC1851_counterAddrOne_13 = (CICC1851_counterAddrOne_14 / 2'b10);
  assign CICC1851_counterAddrOne_14 = ({1'b0,outPixelAddr_value} + CICC1851_counterAddrOne_15);
  assign CICC1851_counterAddrOne_16 = {1'b0,1'b1};
  assign CICC1851_counterAddrOne_15 = {10'd0, CICC1851_counterAddrOne_16};
  assign CICC1851_mainAddrTwo_14 = (CICC1851_mainAddrTwo_15 / 2'b10);
  assign CICC1851_mainAddrTwo_15 = (outPixelAddr_value - 11'h001);
  assign CICC1851_counterAddrOne_17 = (CICC1851_counterAddrOne_18 / 2'b10);
  assign CICC1851_counterAddrOne_18 = (outPixelAddr_value - 11'h001);
  assign CICC1851_mainAddrOne_10 = (CICC1851_mainAddrOne_11 / 2'b10);
  assign CICC1851_mainAddrOne_11 = (outPixelAddr_value - 11'h001);
  assign CICC1851_counterAddrTwo_13 = (CICC1851_counterAddrTwo_14 / 2'b10);
  assign CICC1851_counterAddrTwo_14 = (outPixelAddr_value - 11'h001);
  assign CICC1851_mainAddrOne_12 = (CICC1851_mainAddrOne_13 / 2'b10);
  assign CICC1851_mainAddrOne_13 = ({1'b0,outPixelAddr_value} + CICC1851_mainAddrOne_14);
  assign CICC1851_mainAddrOne_15 = {1'b0,1'b1};
  assign CICC1851_mainAddrOne_14 = {10'd0, CICC1851_mainAddrOne_15};
  assign CICC1851_counterAddrTwo_15 = (CICC1851_counterAddrTwo_16 / 2'b10);
  assign CICC1851_counterAddrTwo_16 = ({1'b0,outPixelAddr_value} + CICC1851_counterAddrTwo_17);
  assign CICC1851_counterAddrTwo_18 = {1'b0,1'b1};
  assign CICC1851_counterAddrTwo_17 = {10'd0, CICC1851_counterAddrTwo_18};
  assign CICC1851_when_SuperResolutionPart1_l664 = {1'd0, outPixelAddr_value};
  assign CICC1851_when_SuperResolutionPart1_l664_1 = (CICC1851_when_SuperResolutionPart1_l664_2 - 12'h002);
  assign CICC1851_when_SuperResolutionPart1_l664_2 = (2'b10 * bmpWidth);
  assign CICC1851_when_SuperResolutionPart1_l665 = {1'd0, outRowCount_value};
  assign CICC1851_when_SuperResolutionPart1_l665_1 = (CICC1851_when_SuperResolutionPart1_l665_2 - 12'h002);
  assign CICC1851_when_SuperResolutionPart1_l665_2 = (2'b10 * bmpHeight);
  assign CICC1851_lineBufferOne_port = passPixels_payload_pixel;
  assign CICC1851_lineBufferOne_port_1 = (passPixels_fire_7 && (! bufferSwitch));
  assign CICC1851_lineBufferTwo_port = passPixels_payload_pixel;
  assign CICC1851_lineBufferTwo_port_1 = (passPixels_fire_6 && bufferSwitch);
  always @(posedge clk) begin
    if(mainAddrOneStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferOne_port0 <= lineBufferOne[mainAddrOneStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(counterAddrOneStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferOne_port1 <= lineBufferOne[counterAddrOneStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(CICC1851_lineBufferOne_port_1) begin
      lineBufferOne[bufferWAddr_value] <= CICC1851_lineBufferOne_port;
    end
  end

  always @(posedge clk) begin
    if(mainAddrTwoStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferTwo_port0 <= lineBufferTwo[mainAddrTwoStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(counterAddrTwoStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferTwo_port1 <= lineBufferTwo[counterAddrTwoStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(CICC1851_lineBufferTwo_port_1) begin
      lineBufferTwo[bufferWAddr_value] <= CICC1851_lineBufferTwo_port;
    end
  end

  StreamFork_1 diffStage_controlPipe_fork (
    .io_input_valid                      (diffStage_controlPipe_valid                                     ), //i
    .io_input_ready                      (diffStage_controlPipe_fork_io_input_ready                       ), //o
    .io_input_payload_frameStart         (diffStage_controlPipe_payload_frameStart                        ), //i
    .io_input_payload_rowEnd             (diffStage_controlPipe_payload_rowEnd                            ), //i
    .io_input_payload_passMode           (diffStage_controlPipe_payload_passMode                          ), //i
    .io_input_payload_passValid          (diffStage_controlPipe_payload_passValid                         ), //i
    .io_input_payload_onceMode           (diffStage_controlPipe_payload_onceMode[2:0]                     ), //i
    .io_input_payload_onceValid          (diffStage_controlPipe_payload_onceValid                         ), //i
    .io_input_payload_mainCompare        (diffStage_controlPipe_payload_mainCompare                       ), //i
    .io_input_payload_counterCompare     (diffStage_controlPipe_payload_counterCompare                    ), //i
    .io_input_payload_mainDiff           (diffStage_controlPipe_payload_mainDiff[7:0]                     ), //i
    .io_input_payload_counterDiff        (diffStage_controlPipe_payload_counterDiff[7:0]                  ), //i
    .io_input_payload_twiceCompValid     (diffStage_controlPipe_payload_twiceCompValid                    ), //i
    .io_input_payload_twiceMode          (diffStage_controlPipe_payload_twiceMode[2:0]                    ), //i
    .io_outputs_0_valid                  (diffStage_controlPipe_fork_io_outputs_0_valid                   ), //o
    .io_outputs_0_ready                  (diffStage_controlPipe_fork_io_outputs_0_ready                   ), //i
    .io_outputs_0_payload_frameStart     (diffStage_controlPipe_fork_io_outputs_0_payload_frameStart      ), //o
    .io_outputs_0_payload_rowEnd         (diffStage_controlPipe_fork_io_outputs_0_payload_rowEnd          ), //o
    .io_outputs_0_payload_passMode       (diffStage_controlPipe_fork_io_outputs_0_payload_passMode        ), //o
    .io_outputs_0_payload_passValid      (diffStage_controlPipe_fork_io_outputs_0_payload_passValid       ), //o
    .io_outputs_0_payload_onceMode       (diffStage_controlPipe_fork_io_outputs_0_payload_onceMode[2:0]   ), //o
    .io_outputs_0_payload_onceValid      (diffStage_controlPipe_fork_io_outputs_0_payload_onceValid       ), //o
    .io_outputs_0_payload_mainCompare    (diffStage_controlPipe_fork_io_outputs_0_payload_mainCompare     ), //o
    .io_outputs_0_payload_counterCompare (diffStage_controlPipe_fork_io_outputs_0_payload_counterCompare  ), //o
    .io_outputs_0_payload_mainDiff       (diffStage_controlPipe_fork_io_outputs_0_payload_mainDiff[7:0]   ), //o
    .io_outputs_0_payload_counterDiff    (diffStage_controlPipe_fork_io_outputs_0_payload_counterDiff[7:0]), //o
    .io_outputs_0_payload_twiceCompValid (diffStage_controlPipe_fork_io_outputs_0_payload_twiceCompValid  ), //o
    .io_outputs_0_payload_twiceMode      (diffStage_controlPipe_fork_io_outputs_0_payload_twiceMode[2:0]  ), //o
    .io_outputs_1_valid                  (diffStage_controlPipe_fork_io_outputs_1_valid                   ), //o
    .io_outputs_1_ready                  (resultStage_pixelStream_ready                                   ), //i
    .io_outputs_1_payload_frameStart     (diffStage_controlPipe_fork_io_outputs_1_payload_frameStart      ), //o
    .io_outputs_1_payload_rowEnd         (diffStage_controlPipe_fork_io_outputs_1_payload_rowEnd          ), //o
    .io_outputs_1_payload_passMode       (diffStage_controlPipe_fork_io_outputs_1_payload_passMode        ), //o
    .io_outputs_1_payload_passValid      (diffStage_controlPipe_fork_io_outputs_1_payload_passValid       ), //o
    .io_outputs_1_payload_onceMode       (diffStage_controlPipe_fork_io_outputs_1_payload_onceMode[2:0]   ), //o
    .io_outputs_1_payload_onceValid      (diffStage_controlPipe_fork_io_outputs_1_payload_onceValid       ), //o
    .io_outputs_1_payload_mainCompare    (diffStage_controlPipe_fork_io_outputs_1_payload_mainCompare     ), //o
    .io_outputs_1_payload_counterCompare (diffStage_controlPipe_fork_io_outputs_1_payload_counterCompare  ), //o
    .io_outputs_1_payload_mainDiff       (diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff[7:0]   ), //o
    .io_outputs_1_payload_counterDiff    (diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff[7:0]), //o
    .io_outputs_1_payload_twiceCompValid (diffStage_controlPipe_fork_io_outputs_1_payload_twiceCompValid  ), //o
    .io_outputs_1_payload_twiceMode      (diffStage_controlPipe_fork_io_outputs_1_payload_twiceMode[2:0]  )  //o
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_3_BOOT : controlStateMachine_stateReg_string = "BOOT ";
      controlStateMachine_enumDef_3_HOLD : controlStateMachine_stateReg_string = "HOLD ";
      controlStateMachine_enumDef_3_PASS : controlStateMachine_stateReg_string = "PASS ";
      controlStateMachine_enumDef_3_ONCE : controlStateMachine_stateReg_string = "ONCE ";
      controlStateMachine_enumDef_3_TWICE : controlStateMachine_stateReg_string = "TWICE";
      default : controlStateMachine_stateReg_string = "?????";
    endcase
  end
  always @(*) begin
    case(controlStateMachine_stateNext)
      controlStateMachine_enumDef_3_BOOT : controlStateMachine_stateNext_string = "BOOT ";
      controlStateMachine_enumDef_3_HOLD : controlStateMachine_stateNext_string = "HOLD ";
      controlStateMachine_enumDef_3_PASS : controlStateMachine_stateNext_string = "PASS ";
      controlStateMachine_enumDef_3_ONCE : controlStateMachine_stateNext_string = "ONCE ";
      controlStateMachine_enumDef_3_TWICE : controlStateMachine_stateNext_string = "TWICE";
      default : controlStateMachine_stateNext_string = "?????";
    endcase
  end
  `endif

  always @(*) begin
    pixelsIn_ready = 1'b0;
    pixelsIn_ready = (! pixelsIn_rValid);
  end

  always @(*) begin
    pixelsOut_valid = 1'b0;
    pixelsOut_valid = pixelsStream_s2mPipe_m2sPipe_valid;
  end

  always @(*) begin
    pixelsOut_payload_pixel = 8'h0;
    pixelsOut_payload_pixel = pixelsStream_s2mPipe_m2sPipe_payload_pixel;
  end

  always @(*) begin
    pixelsOut_payload_frameStart = 1'b0;
    pixelsOut_payload_frameStart = pixelsStream_s2mPipe_m2sPipe_payload_frameStart;
  end

  always @(*) begin
    pixelsOut_payload_rowEnd = 1'b0;
    pixelsOut_payload_rowEnd = pixelsStream_s2mPipe_m2sPipe_payload_rowEnd;
  end

  always @(*) begin
    startOut = 1'b0;
    startOut = slaveStart;
  end

  always @(*) begin
    inpDoneOut = 1'b0;
    inpDoneOut = inpDone;
  end

  assign when_SuperResolutionPart1_l79 = (inpThreeDoneIn && inpTwoDoneIn);
  assign when_SuperResolutionPart1_l79_1 = (startIn && (! startIn_regNext));
  assign when_SuperResolutionPart1_l82 = (! startIn);
  assign when_SuperResolutionPart1_l85 = (startIn && (! readDone));
  assign when_SuperResolutionPart1_l85_1 = (! startIn);
  assign pixelsIn_fire = (pixelsIn_valid && pixelsIn_ready);
  assign when_SuperResolutionPart1_l88 = ((! inpTwoDoneIn) && pixelsIn_fire);
  assign when_SuperResolutionPart1_l88_1 = ((inpTwoDoneIn && inpThreeDoneIn) || (! startIn));
  assign when_SuperResolutionPart1_l103 = (! startIn);
  assign when_SuperResolutionPart1_l106 = (! startIn);
  always @(*) begin
    bufferRowCount_willIncrement = 1'b0;
    if(when_SuperResolutionPart1_l425) begin
      if(!bufferReachFinalRow) begin
        bufferRowCount_willIncrement = 1'b1;
      end
    end
  end

  always @(*) begin
    bufferRowCount_willClear = 1'b0;
    if(when_SuperResolutionPart1_l425) begin
      if(bufferReachFinalRow) begin
        bufferRowCount_willClear = 1'b1;
      end
    end
  end

  assign bufferRowCount_willOverflowIfInc = (bufferRowCount_value == 10'h21c);
  assign bufferRowCount_willOverflow = (bufferRowCount_willOverflowIfInc && bufferRowCount_willIncrement);
  always @(*) begin
    if(bufferRowCount_willOverflow) begin
      bufferRowCount_valueNext = 10'h0;
    end else begin
      bufferRowCount_valueNext = (bufferRowCount_value + CICC1851_bufferRowCount_valueNext);
    end
    if(bufferRowCount_willClear) begin
      bufferRowCount_valueNext = 10'h0;
    end
  end

  assign when_SuperResolutionPart1_l112 = ((startIn && (! holdBuffer)) && (! writeDone));
  assign when_SuperResolutionPart1_l112_1 = (((! startIn) || holdBuffer) || writeDone);
  assign when_SuperResolutionPart1_l115 = (! startRead);
  assign when_SuperResolutionPart1_l118 = (! startRead);
  always @(*) begin
    bufferWAddr_willIncrement = 1'b0;
    if(passPixels_fire_8) begin
      if(!passPixels_payload_rowEnd) begin
        bufferWAddr_willIncrement = 1'b1;
      end
    end
  end

  always @(*) begin
    bufferWAddr_willClear = 1'b0;
    if(passPixels_fire_8) begin
      if(passPixels_payload_rowEnd) begin
        bufferWAddr_willClear = 1'b1;
      end
    end
  end

  assign bufferWAddr_willOverflowIfInc = (bufferWAddr_value == 10'h3bf);
  assign bufferWAddr_willOverflow = (bufferWAddr_willOverflowIfInc && bufferWAddr_willIncrement);
  always @(*) begin
    if(bufferWAddr_willOverflow) begin
      bufferWAddr_valueNext = 10'h0;
    end else begin
      bufferWAddr_valueNext = (bufferWAddr_value + CICC1851_bufferWAddr_valueNext);
    end
    if(bufferWAddr_willClear) begin
      bufferWAddr_valueNext = 10'h0;
    end
  end

  always @(*) begin
    outPixelAddr_willIncrement = 1'b0;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_3_HOLD : begin
      end
      controlStateMachine_enumDef_3_PASS : begin
        if(controlStream_fire_6) begin
          if(!outReachRowEnd) begin
            outPixelAddr_willIncrement = 1'b1;
          end
        end
      end
      controlStateMachine_enumDef_3_ONCE : begin
        if(controlStream_fire_12) begin
          if(!outReachRowEnd) begin
            outPixelAddr_willIncrement = 1'b1;
          end
        end
      end
      controlStateMachine_enumDef_3_TWICE : begin
        if(controlStream_fire_17) begin
          if(!outReachRowEnd) begin
            outPixelAddr_willIncrement = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outPixelAddr_willClear = 1'b0;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_3_HOLD : begin
      end
      controlStateMachine_enumDef_3_PASS : begin
        if(controlStream_fire_6) begin
          if(outReachRowEnd) begin
            outPixelAddr_willClear = 1'b1;
          end
        end
      end
      controlStateMachine_enumDef_3_ONCE : begin
        if(controlStream_fire_12) begin
          if(outReachRowEnd) begin
            outPixelAddr_willClear = 1'b1;
          end
        end
      end
      controlStateMachine_enumDef_3_TWICE : begin
        if(controlStream_fire_17) begin
          if(outReachRowEnd) begin
            outPixelAddr_willClear = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign outPixelAddr_willOverflowIfInc = (outPixelAddr_value == 11'h77f);
  assign outPixelAddr_willOverflow = (outPixelAddr_willOverflowIfInc && outPixelAddr_willIncrement);
  always @(*) begin
    if(outPixelAddr_willOverflow) begin
      outPixelAddr_valueNext = 11'h0;
    end else begin
      outPixelAddr_valueNext = (outPixelAddr_value + CICC1851_outPixelAddr_valueNext);
    end
    if(outPixelAddr_willClear) begin
      outPixelAddr_valueNext = 11'h0;
    end
  end

  always @(*) begin
    outRowCount_willIncrement = 1'b0;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_3_HOLD : begin
      end
      controlStateMachine_enumDef_3_PASS : begin
        if(when_SuperResolutionPart1_l513) begin
          if(!outReachFinalRow) begin
            outRowCount_willIncrement = 1'b1;
          end
        end
      end
      controlStateMachine_enumDef_3_ONCE : begin
        if(when_SuperResolutionPart1_l581) begin
          if(!outReachFinalRow) begin
            outRowCount_willIncrement = 1'b1;
          end
        end
      end
      controlStateMachine_enumDef_3_TWICE : begin
        if(when_SuperResolutionPart1_l667) begin
          if(!outReachFinalRow) begin
            outRowCount_willIncrement = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outRowCount_willClear = 1'b0;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_3_HOLD : begin
      end
      controlStateMachine_enumDef_3_PASS : begin
        if(when_SuperResolutionPart1_l513) begin
          if(outReachFinalRow) begin
            outRowCount_willClear = 1'b1;
          end
        end
      end
      controlStateMachine_enumDef_3_ONCE : begin
        if(when_SuperResolutionPart1_l581) begin
          if(outReachFinalRow) begin
            outRowCount_willClear = 1'b1;
          end
        end
      end
      controlStateMachine_enumDef_3_TWICE : begin
        if(when_SuperResolutionPart1_l667) begin
          if(outReachFinalRow) begin
            outRowCount_willClear = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign outRowCount_willOverflowIfInc = (outRowCount_value == 11'h438);
  assign outRowCount_willOverflow = (outRowCount_willOverflowIfInc && outRowCount_willIncrement);
  always @(*) begin
    if(outRowCount_willOverflow) begin
      outRowCount_valueNext = 11'h0;
    end else begin
      outRowCount_valueNext = (outRowCount_value + CICC1851_outRowCount_valueNext);
    end
    if(outRowCount_willClear) begin
      outRowCount_valueNext = 11'h0;
    end
  end

  always @(*) begin
    mainAddrOne = CICC1851_mainAddrOne[9:0];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_3_HOLD : begin
      end
      controlStateMachine_enumDef_3_PASS : begin
      end
      controlStateMachine_enumDef_3_ONCE : begin
        if(when_SuperResolutionPart1_l537) begin
          if(nextRowBuffer) begin
            mainAddrOne = CICC1851_mainAddrOne_1[9:0];
          end
        end else begin
          mainAddrOne = CICC1851_mainAddrOne_3[9:0];
        end
      end
      controlStateMachine_enumDef_3_TWICE : begin
        if(outReachFinalRow) begin
          if(nextRowBuffer) begin
            if(outReachRowEnd) begin
              mainAddrOne = CICC1851_mainAddrOne_4[9:0];
            end else begin
              mainAddrOne = CICC1851_mainAddrOne_6[9:0];
            end
          end
        end else begin
          if(nextRowBuffer) begin
            mainAddrOne = CICC1851_mainAddrOne_8[9:0];
          end else begin
            if(outReachRowEnd) begin
              mainAddrOne = CICC1851_mainAddrOne_10[9:0];
            end else begin
              mainAddrOne = CICC1851_mainAddrOne_12[9:0];
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    counterAddrOne = CICC1851_counterAddrOne[9:0];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_3_HOLD : begin
      end
      controlStateMachine_enumDef_3_PASS : begin
      end
      controlStateMachine_enumDef_3_ONCE : begin
        if(when_SuperResolutionPart1_l537) begin
          if(nextRowBuffer) begin
            if(outReachRowEnd) begin
              counterAddrOne = CICC1851_counterAddrOne_1[9:0];
            end else begin
              counterAddrOne = CICC1851_counterAddrOne_3[9:0];
            end
          end
        end
      end
      controlStateMachine_enumDef_3_TWICE : begin
        if(outReachFinalRow) begin
          if(nextRowBuffer) begin
            if(!outReachRowEnd) begin
              counterAddrOne = CICC1851_counterAddrOne_7[9:0];
            end
          end
        end else begin
          if(nextRowBuffer) begin
            if(outReachRowEnd) begin
              counterAddrOne = CICC1851_counterAddrOne_11[9:0];
            end else begin
              counterAddrOne = CICC1851_counterAddrOne_13[9:0];
            end
          end else begin
            counterAddrOne = CICC1851_counterAddrOne_17[9:0];
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    mainAddrTwo = CICC1851_mainAddrTwo[9:0];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_3_HOLD : begin
      end
      controlStateMachine_enumDef_3_PASS : begin
      end
      controlStateMachine_enumDef_3_ONCE : begin
        if(when_SuperResolutionPart1_l537) begin
          if(!nextRowBuffer) begin
            mainAddrTwo = CICC1851_mainAddrTwo_1[9:0];
          end
        end else begin
          mainAddrTwo = CICC1851_mainAddrTwo_3[9:0];
        end
      end
      controlStateMachine_enumDef_3_TWICE : begin
        if(outReachFinalRow) begin
          if(!nextRowBuffer) begin
            if(outReachRowEnd) begin
              mainAddrTwo = CICC1851_mainAddrTwo_4[9:0];
            end else begin
              mainAddrTwo = CICC1851_mainAddrTwo_6[9:0];
            end
          end
        end else begin
          if(nextRowBuffer) begin
            if(outReachRowEnd) begin
              mainAddrTwo = CICC1851_mainAddrTwo_8[9:0];
            end else begin
              mainAddrTwo = CICC1851_mainAddrTwo_10[9:0];
            end
          end else begin
            mainAddrTwo = CICC1851_mainAddrTwo_14[9:0];
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    counterAddrTwo = CICC1851_counterAddrTwo[9:0];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_3_HOLD : begin
      end
      controlStateMachine_enumDef_3_PASS : begin
      end
      controlStateMachine_enumDef_3_ONCE : begin
        if(when_SuperResolutionPart1_l537) begin
          if(!nextRowBuffer) begin
            if(outReachRowEnd) begin
              counterAddrTwo = CICC1851_counterAddrTwo_1[9:0];
            end else begin
              counterAddrTwo = CICC1851_counterAddrTwo_3[9:0];
            end
          end
        end
      end
      controlStateMachine_enumDef_3_TWICE : begin
        if(outReachFinalRow) begin
          if(!nextRowBuffer) begin
            if(!outReachRowEnd) begin
              counterAddrTwo = CICC1851_counterAddrTwo_7[9:0];
            end
          end
        end else begin
          if(nextRowBuffer) begin
            counterAddrTwo = CICC1851_counterAddrTwo_11[9:0];
          end else begin
            if(outReachRowEnd) begin
              counterAddrTwo = CICC1851_counterAddrTwo_13[9:0];
            end else begin
              counterAddrTwo = CICC1851_counterAddrTwo_15[9:0];
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign validStream_valid = 1'b1;
  assign CICC1851_controls_frameStart = 30'h0;
  always @(*) begin
    controls_frameStart = CICC1851_controls_frameStart[0];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_3_HOLD : begin
      end
      controlStateMachine_enumDef_3_PASS : begin
        if(frameStart) begin
          controls_frameStart = 1'b1;
        end
      end
      controlStateMachine_enumDef_3_ONCE : begin
      end
      controlStateMachine_enumDef_3_TWICE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_rowEnd = CICC1851_controls_frameStart[1];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_3_HOLD : begin
      end
      controlStateMachine_enumDef_3_PASS : begin
        if(outReachRowEnd) begin
          controls_rowEnd = 1'b1;
        end
      end
      controlStateMachine_enumDef_3_ONCE : begin
        if(outReachRowEnd) begin
          controls_rowEnd = 1'b1;
        end
      end
      controlStateMachine_enumDef_3_TWICE : begin
        if(outReachRowEnd) begin
          controls_rowEnd = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_passMode = CICC1851_controls_frameStart[2];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_3_HOLD : begin
      end
      controlStateMachine_enumDef_3_PASS : begin
        if(nextRowBuffer) begin
          controls_passMode = 1'b0;
        end else begin
          controls_passMode = 1'b1;
        end
      end
      controlStateMachine_enumDef_3_ONCE : begin
      end
      controlStateMachine_enumDef_3_TWICE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_passValid = CICC1851_controls_frameStart[3];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_3_HOLD : begin
      end
      controlStateMachine_enumDef_3_PASS : begin
        controls_passValid = 1'b1;
      end
      controlStateMachine_enumDef_3_ONCE : begin
      end
      controlStateMachine_enumDef_3_TWICE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_onceMode = CICC1851_controls_frameStart[6 : 4];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_3_HOLD : begin
      end
      controlStateMachine_enumDef_3_PASS : begin
      end
      controlStateMachine_enumDef_3_ONCE : begin
        if(when_SuperResolutionPart1_l537) begin
          if(nextRowBuffer) begin
            controls_onceMode = 3'b000;
          end else begin
            controls_onceMode = {2'd0, CICC1851_controls_onceMode};
          end
        end else begin
          if(outReachFinalRow) begin
            if(nextRowBuffer) begin
              controls_onceMode = 3'b101;
            end else begin
              controls_onceMode = 3'b100;
            end
          end else begin
            if(nextRowBuffer) begin
              controls_onceMode = {1'd0, CICC1851_controls_onceMode_1};
            end else begin
              controls_onceMode = {1'd0, CICC1851_controls_onceMode_2};
            end
          end
        end
      end
      controlStateMachine_enumDef_3_TWICE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_onceValid = CICC1851_controls_frameStart[7];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_3_HOLD : begin
      end
      controlStateMachine_enumDef_3_PASS : begin
      end
      controlStateMachine_enumDef_3_ONCE : begin
        controls_onceValid = 1'b1;
      end
      controlStateMachine_enumDef_3_TWICE : begin
      end
      default : begin
      end
    endcase
  end

  assign controls_mainCompare = CICC1851_controls_frameStart[8];
  assign controls_counterCompare = CICC1851_controls_frameStart[9];
  assign controls_mainDiff = CICC1851_controls_frameStart[17 : 10];
  assign controls_counterDiff = CICC1851_controls_frameStart[25 : 18];
  always @(*) begin
    controls_twiceCompValid = CICC1851_controls_frameStart[26];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_3_HOLD : begin
      end
      controlStateMachine_enumDef_3_PASS : begin
      end
      controlStateMachine_enumDef_3_ONCE : begin
      end
      controlStateMachine_enumDef_3_TWICE : begin
        controls_twiceCompValid = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_twiceMode = CICC1851_controls_frameStart[29 : 27];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_3_HOLD : begin
      end
      controlStateMachine_enumDef_3_PASS : begin
      end
      controlStateMachine_enumDef_3_ONCE : begin
      end
      controlStateMachine_enumDef_3_TWICE : begin
        if(outReachFinalRow) begin
          if(nextRowBuffer) begin
            if(outReachRowEnd) begin
              controls_twiceMode = 3'b100;
            end else begin
              controls_twiceMode = 3'b101;
            end
          end else begin
            if(outReachRowEnd) begin
              controls_twiceMode = 3'b010;
            end else begin
              controls_twiceMode = 3'b011;
            end
          end
        end else begin
          if(nextRowBuffer) begin
            controls_twiceMode = 3'b000;
          end else begin
            controls_twiceMode = 3'b001;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    validStream_ready = (controlStream_ready && startRead);
    validStream_ready = (mainAddrOneStream_ready && startRead);
    validStream_ready = (counterAddrOneStream_ready && startRead);
    validStream_ready = (mainAddrTwoStream_ready && startRead);
    validStream_ready = (counterAddrTwoStream_ready && startRead);
  end

  assign controlStream_valid = (validStream_valid && startRead);
  assign controlStream_payload_frameStart = controls_frameStart;
  assign controlStream_payload_rowEnd = controls_rowEnd;
  assign controlStream_payload_passMode = controls_passMode;
  assign controlStream_payload_passValid = controls_passValid;
  assign controlStream_payload_onceMode = controls_onceMode;
  assign controlStream_payload_onceValid = controls_onceValid;
  assign controlStream_payload_mainCompare = controls_mainCompare;
  assign controlStream_payload_counterCompare = controls_counterCompare;
  assign controlStream_payload_mainDiff = controls_mainDiff;
  assign controlStream_payload_counterDiff = controls_counterDiff;
  assign controlStream_payload_twiceCompValid = controls_twiceCompValid;
  assign controlStream_payload_twiceMode = controls_twiceMode;
  assign mainAddrOneStream_valid = (validStream_valid && startRead);
  assign mainAddrOneStream_payload = mainAddrOne;
  assign counterAddrOneStream_valid = (validStream_valid && startRead);
  assign counterAddrOneStream_payload = counterAddrOne;
  assign mainAddrTwoStream_valid = (validStream_valid && startRead);
  assign mainAddrTwoStream_payload = mainAddrTwo;
  assign counterAddrTwoStream_valid = (validStream_valid && startRead);
  assign counterAddrTwoStream_payload = counterAddrTwo;
  assign mainAddrOneStream_ready = (! mainAddrOneStream_rValid);
  assign mainAddrOneStream_s2mPipe_valid = (mainAddrOneStream_valid || mainAddrOneStream_rValid);
  assign mainAddrOneStream_s2mPipe_payload = (mainAddrOneStream_rValid ? mainAddrOneStream_rData : mainAddrOneStream_payload);
  always @(*) begin
    mainAddrOneStream_s2mPipe_ready = mainAddrOneStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368) begin
      mainAddrOneStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368 = (! mainAddrOneStream_s2mPipe_m2sPipe_valid);
  assign mainAddrOneStream_s2mPipe_m2sPipe_valid = mainAddrOneStream_s2mPipe_rValid;
  assign mainAddrOneStream_s2mPipe_m2sPipe_payload = mainAddrOneStream_s2mPipe_rData;
  assign mainAddrOneStream_s2mPipe_m2sPipe_ready = ((! CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready) || CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready = CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_mainOnePixelStream_payload = CICC1851_lineBufferOne_port0;
  assign CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_1 = readStage_mainOnePixelStream_ready;
    if(when_Stream_l368_1) begin
      CICC1851_1 = 1'b1;
    end
  end

  assign when_Stream_l368_1 = (! readStage_mainOnePixelStream_valid);
  assign readStage_mainOnePixelStream_valid = CICC1851_readStage_mainOnePixelStream_valid;
  assign readStage_mainOnePixelStream_payload = CICC1851_readStage_mainOnePixelStream_payload_2;
  assign counterAddrOneStream_ready = (! counterAddrOneStream_rValid);
  assign counterAddrOneStream_s2mPipe_valid = (counterAddrOneStream_valid || counterAddrOneStream_rValid);
  assign counterAddrOneStream_s2mPipe_payload = (counterAddrOneStream_rValid ? counterAddrOneStream_rData : counterAddrOneStream_payload);
  always @(*) begin
    counterAddrOneStream_s2mPipe_ready = counterAddrOneStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_2) begin
      counterAddrOneStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_2 = (! counterAddrOneStream_s2mPipe_m2sPipe_valid);
  assign counterAddrOneStream_s2mPipe_m2sPipe_valid = counterAddrOneStream_s2mPipe_rValid;
  assign counterAddrOneStream_s2mPipe_m2sPipe_payload = counterAddrOneStream_s2mPipe_rData;
  assign counterAddrOneStream_s2mPipe_m2sPipe_ready = ((! CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready) || CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready = CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_counterOnePixelStream_payload = CICC1851_lineBufferOne_port1;
  assign CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_2 = readStage_counterOnePixelStream_ready;
    if(when_Stream_l368_3) begin
      CICC1851_2 = 1'b1;
    end
  end

  assign when_Stream_l368_3 = (! readStage_counterOnePixelStream_valid);
  assign readStage_counterOnePixelStream_valid = CICC1851_readStage_counterOnePixelStream_valid;
  assign readStage_counterOnePixelStream_payload = CICC1851_readStage_counterOnePixelStream_payload_2;
  assign mainAddrTwoStream_ready = (! mainAddrTwoStream_rValid);
  assign mainAddrTwoStream_s2mPipe_valid = (mainAddrTwoStream_valid || mainAddrTwoStream_rValid);
  assign mainAddrTwoStream_s2mPipe_payload = (mainAddrTwoStream_rValid ? mainAddrTwoStream_rData : mainAddrTwoStream_payload);
  always @(*) begin
    mainAddrTwoStream_s2mPipe_ready = mainAddrTwoStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_4) begin
      mainAddrTwoStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_4 = (! mainAddrTwoStream_s2mPipe_m2sPipe_valid);
  assign mainAddrTwoStream_s2mPipe_m2sPipe_valid = mainAddrTwoStream_s2mPipe_rValid;
  assign mainAddrTwoStream_s2mPipe_m2sPipe_payload = mainAddrTwoStream_s2mPipe_rData;
  assign mainAddrTwoStream_s2mPipe_m2sPipe_ready = ((! CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready) || CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready = CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_mainTwoPixelStream_payload = CICC1851_lineBufferTwo_port0;
  assign CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_3 = readStage_mainTwoPixelStream_ready;
    if(when_Stream_l368_5) begin
      CICC1851_3 = 1'b1;
    end
  end

  assign when_Stream_l368_5 = (! readStage_mainTwoPixelStream_valid);
  assign readStage_mainTwoPixelStream_valid = CICC1851_readStage_mainTwoPixelStream_valid;
  assign readStage_mainTwoPixelStream_payload = CICC1851_readStage_mainTwoPixelStream_payload_2;
  assign counterAddrTwoStream_ready = (! counterAddrTwoStream_rValid);
  assign counterAddrTwoStream_s2mPipe_valid = (counterAddrTwoStream_valid || counterAddrTwoStream_rValid);
  assign counterAddrTwoStream_s2mPipe_payload = (counterAddrTwoStream_rValid ? counterAddrTwoStream_rData : counterAddrTwoStream_payload);
  always @(*) begin
    counterAddrTwoStream_s2mPipe_ready = counterAddrTwoStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_6) begin
      counterAddrTwoStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_6 = (! counterAddrTwoStream_s2mPipe_m2sPipe_valid);
  assign counterAddrTwoStream_s2mPipe_m2sPipe_valid = counterAddrTwoStream_s2mPipe_rValid;
  assign counterAddrTwoStream_s2mPipe_m2sPipe_payload = counterAddrTwoStream_s2mPipe_rData;
  assign counterAddrTwoStream_s2mPipe_m2sPipe_ready = ((! CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready) || CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready = CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_counterTwoPixelStream_payload = CICC1851_lineBufferTwo_port1;
  assign CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_4 = readStage_counterTwoPixelStream_ready;
    if(when_Stream_l368_7) begin
      CICC1851_4 = 1'b1;
    end
  end

  assign when_Stream_l368_7 = (! readStage_counterTwoPixelStream_valid);
  assign readStage_counterTwoPixelStream_valid = CICC1851_readStage_counterTwoPixelStream_valid;
  assign readStage_counterTwoPixelStream_payload = CICC1851_readStage_counterTwoPixelStream_payload_2;
  assign controlStream_ready = (! controlStream_rValid);
  assign controlStream_s2mPipe_valid = (controlStream_valid || controlStream_rValid);
  assign controlStream_s2mPipe_payload_frameStart = (controlStream_rValid ? controlStream_rData_frameStart : controlStream_payload_frameStart);
  assign controlStream_s2mPipe_payload_rowEnd = (controlStream_rValid ? controlStream_rData_rowEnd : controlStream_payload_rowEnd);
  assign controlStream_s2mPipe_payload_passMode = (controlStream_rValid ? controlStream_rData_passMode : controlStream_payload_passMode);
  assign controlStream_s2mPipe_payload_passValid = (controlStream_rValid ? controlStream_rData_passValid : controlStream_payload_passValid);
  assign controlStream_s2mPipe_payload_onceMode = (controlStream_rValid ? controlStream_rData_onceMode : controlStream_payload_onceMode);
  assign controlStream_s2mPipe_payload_onceValid = (controlStream_rValid ? controlStream_rData_onceValid : controlStream_payload_onceValid);
  assign controlStream_s2mPipe_payload_mainCompare = (controlStream_rValid ? controlStream_rData_mainCompare : controlStream_payload_mainCompare);
  assign controlStream_s2mPipe_payload_counterCompare = (controlStream_rValid ? controlStream_rData_counterCompare : controlStream_payload_counterCompare);
  assign controlStream_s2mPipe_payload_mainDiff = (controlStream_rValid ? controlStream_rData_mainDiff : controlStream_payload_mainDiff);
  assign controlStream_s2mPipe_payload_counterDiff = (controlStream_rValid ? controlStream_rData_counterDiff : controlStream_payload_counterDiff);
  assign controlStream_s2mPipe_payload_twiceCompValid = (controlStream_rValid ? controlStream_rData_twiceCompValid : controlStream_payload_twiceCompValid);
  assign controlStream_s2mPipe_payload_twiceMode = (controlStream_rValid ? controlStream_rData_twiceMode : controlStream_payload_twiceMode);
  always @(*) begin
    controlStream_s2mPipe_ready = controlStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_8) begin
      controlStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_8 = (! controlStream_s2mPipe_m2sPipe_valid);
  assign controlStream_s2mPipe_m2sPipe_valid = controlStream_s2mPipe_rValid;
  assign controlStream_s2mPipe_m2sPipe_payload_frameStart = controlStream_s2mPipe_rData_frameStart;
  assign controlStream_s2mPipe_m2sPipe_payload_rowEnd = controlStream_s2mPipe_rData_rowEnd;
  assign controlStream_s2mPipe_m2sPipe_payload_passMode = controlStream_s2mPipe_rData_passMode;
  assign controlStream_s2mPipe_m2sPipe_payload_passValid = controlStream_s2mPipe_rData_passValid;
  assign controlStream_s2mPipe_m2sPipe_payload_onceMode = controlStream_s2mPipe_rData_onceMode;
  assign controlStream_s2mPipe_m2sPipe_payload_onceValid = controlStream_s2mPipe_rData_onceValid;
  assign controlStream_s2mPipe_m2sPipe_payload_mainCompare = controlStream_s2mPipe_rData_mainCompare;
  assign controlStream_s2mPipe_m2sPipe_payload_counterCompare = controlStream_s2mPipe_rData_counterCompare;
  assign controlStream_s2mPipe_m2sPipe_payload_mainDiff = controlStream_s2mPipe_rData_mainDiff;
  assign controlStream_s2mPipe_m2sPipe_payload_counterDiff = controlStream_s2mPipe_rData_counterDiff;
  assign controlStream_s2mPipe_m2sPipe_payload_twiceCompValid = controlStream_s2mPipe_rData_twiceCompValid;
  assign controlStream_s2mPipe_m2sPipe_payload_twiceMode = controlStream_s2mPipe_rData_twiceMode;
  always @(*) begin
    controlStream_s2mPipe_m2sPipe_ready = controlStream_s2mPipe_m2sPipe_m2sPipe_ready;
    if(when_Stream_l368_9) begin
      controlStream_s2mPipe_m2sPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_9 = (! controlStream_s2mPipe_m2sPipe_m2sPipe_valid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_valid = controlStream_s2mPipe_m2sPipe_rValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_frameStart = controlStream_s2mPipe_m2sPipe_rData_frameStart;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_rowEnd = controlStream_s2mPipe_m2sPipe_rData_rowEnd;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passMode = controlStream_s2mPipe_m2sPipe_rData_passMode;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passValid = controlStream_s2mPipe_m2sPipe_rData_passValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceMode = controlStream_s2mPipe_m2sPipe_rData_onceMode;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceValid = controlStream_s2mPipe_m2sPipe_rData_onceValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainCompare = controlStream_s2mPipe_m2sPipe_rData_mainCompare;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterCompare = controlStream_s2mPipe_m2sPipe_rData_counterCompare;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDiff = controlStream_s2mPipe_m2sPipe_rData_mainDiff;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDiff = controlStream_s2mPipe_m2sPipe_rData_counterDiff;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceCompValid = controlStream_s2mPipe_m2sPipe_rData_twiceCompValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceMode = controlStream_s2mPipe_m2sPipe_rData_twiceMode;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_ready = (! controlStream_s2mPipe_m2sPipe_m2sPipe_rValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_valid = (controlStream_s2mPipe_m2sPipe_m2sPipe_valid || controlStream_s2mPipe_m2sPipe_m2sPipe_rValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_frameStart = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_frameStart : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_frameStart);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_rowEnd = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_rowEnd : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_rowEnd);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_passMode = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_passMode : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passMode);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_passValid = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_passValid : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_onceMode = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_onceMode : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceMode);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_onceValid = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_onceValid : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainCompare = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainCompare : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainCompare);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterCompare = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterCompare : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterCompare);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainDiff = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainDiff : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDiff);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterDiff = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterDiff : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDiff);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_twiceCompValid = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_twiceCompValid : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceCompValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_twiceMode = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_twiceMode : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceMode);
  always @(*) begin
    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready = readStage_controlPipe_ready;
    if(when_Stream_l368_10) begin
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_10 = (! readStage_controlPipe_valid);
  assign readStage_controlPipe_valid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rValid;
  assign readStage_controlPipe_payload_frameStart = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_frameStart;
  assign readStage_controlPipe_payload_rowEnd = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_rowEnd;
  assign readStage_controlPipe_payload_passMode = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_passMode;
  assign readStage_controlPipe_payload_passValid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_passValid;
  assign readStage_controlPipe_payload_onceMode = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_onceMode;
  assign readStage_controlPipe_payload_onceValid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_onceValid;
  assign readStage_controlPipe_payload_mainCompare = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainCompare;
  assign readStage_controlPipe_payload_counterCompare = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterCompare;
  assign readStage_controlPipe_payload_mainDiff = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainDiff;
  assign readStage_controlPipe_payload_counterDiff = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterDiff;
  assign readStage_controlPipe_payload_twiceCompValid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_twiceCompValid;
  assign readStage_controlPipe_payload_twiceMode = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_twiceMode;
  assign readStage_mainOnePixelStream_ready = (! readStage_mainOnePixelStream_rValid);
  assign readStage_mainOnePixelStream_s2mPipe_valid = (readStage_mainOnePixelStream_valid || readStage_mainOnePixelStream_rValid);
  assign readStage_mainOnePixelStream_s2mPipe_payload = (readStage_mainOnePixelStream_rValid ? readStage_mainOnePixelStream_rData : readStage_mainOnePixelStream_payload);
  always @(*) begin
    readStage_mainOnePixelStream_s2mPipe_ready = compareStage_mainOnePixelStream_ready;
    if(when_Stream_l368_11) begin
      readStage_mainOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_11 = (! compareStage_mainOnePixelStream_valid);
  assign compareStage_mainOnePixelStream_valid = readStage_mainOnePixelStream_s2mPipe_rValid;
  assign compareStage_mainOnePixelStream_payload = readStage_mainOnePixelStream_s2mPipe_rData;
  assign readStage_counterOnePixelStream_ready = (! readStage_counterOnePixelStream_rValid);
  assign readStage_counterOnePixelStream_s2mPipe_valid = (readStage_counterOnePixelStream_valid || readStage_counterOnePixelStream_rValid);
  assign readStage_counterOnePixelStream_s2mPipe_payload = (readStage_counterOnePixelStream_rValid ? readStage_counterOnePixelStream_rData : readStage_counterOnePixelStream_payload);
  always @(*) begin
    readStage_counterOnePixelStream_s2mPipe_ready = compareStage_counterOnePixelStream_ready;
    if(when_Stream_l368_12) begin
      readStage_counterOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_12 = (! compareStage_counterOnePixelStream_valid);
  assign compareStage_counterOnePixelStream_valid = readStage_counterOnePixelStream_s2mPipe_rValid;
  assign compareStage_counterOnePixelStream_payload = readStage_counterOnePixelStream_s2mPipe_rData;
  assign readStage_mainTwoPixelStream_ready = (! readStage_mainTwoPixelStream_rValid);
  assign readStage_mainTwoPixelStream_s2mPipe_valid = (readStage_mainTwoPixelStream_valid || readStage_mainTwoPixelStream_rValid);
  assign readStage_mainTwoPixelStream_s2mPipe_payload = (readStage_mainTwoPixelStream_rValid ? readStage_mainTwoPixelStream_rData : readStage_mainTwoPixelStream_payload);
  always @(*) begin
    readStage_mainTwoPixelStream_s2mPipe_ready = compareStage_mainTwoPixelStream_ready;
    if(when_Stream_l368_13) begin
      readStage_mainTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_13 = (! compareStage_mainTwoPixelStream_valid);
  assign compareStage_mainTwoPixelStream_valid = readStage_mainTwoPixelStream_s2mPipe_rValid;
  assign compareStage_mainTwoPixelStream_payload = readStage_mainTwoPixelStream_s2mPipe_rData;
  assign readStage_counterTwoPixelStream_ready = (! readStage_counterTwoPixelStream_rValid);
  assign readStage_counterTwoPixelStream_s2mPipe_valid = (readStage_counterTwoPixelStream_valid || readStage_counterTwoPixelStream_rValid);
  assign readStage_counterTwoPixelStream_s2mPipe_payload = (readStage_counterTwoPixelStream_rValid ? readStage_counterTwoPixelStream_rData : readStage_counterTwoPixelStream_payload);
  always @(*) begin
    readStage_counterTwoPixelStream_s2mPipe_ready = compareStage_counterTwoPixelStream_ready;
    if(when_Stream_l368_14) begin
      readStage_counterTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_14 = (! compareStage_counterTwoPixelStream_valid);
  assign compareStage_counterTwoPixelStream_valid = readStage_counterTwoPixelStream_s2mPipe_rValid;
  assign compareStage_counterTwoPixelStream_payload = readStage_counterTwoPixelStream_s2mPipe_rData;
  always @(*) begin
    CICC1851_readStage_controlPipe_translated_payload_mainCompare = readStage_controlPipe_payload_mainCompare;
    if(readStage_controlPipe_payload_onceValid) begin
      case(readStage_controlPipe_payload_onceMode)
        3'b000 : begin
          if(when_SuperResolutionPart1_l205) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        3'b001 : begin
          if(when_SuperResolutionPart1_l209) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        3'b010 : begin
          if(when_SuperResolutionPart1_l213) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        3'b011 : begin
          if(when_SuperResolutionPart1_l217) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        3'b100 : begin
          CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
        end
        3'b101 : begin
          CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
        end
        default : begin
        end
      endcase
    end
    if(readStage_controlPipe_payload_twiceCompValid) begin
      case(readStage_controlPipe_payload_twiceMode)
        3'b000 : begin
          if(when_SuperResolutionPart1_l228) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        3'b001 : begin
          if(when_SuperResolutionPart1_l234) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        3'b010 : begin
          CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
        end
        3'b011 : begin
          if(when_SuperResolutionPart1_l241) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        3'b100 : begin
          CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
        end
        3'b101 : begin
          if(when_SuperResolutionPart1_l246) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    CICC1851_readStage_controlPipe_translated_payload_counterCompare = readStage_controlPipe_payload_counterCompare;
    if(readStage_controlPipe_payload_twiceCompValid) begin
      case(readStage_controlPipe_payload_twiceMode)
        3'b000 : begin
          if(when_SuperResolutionPart1_l230) begin
            CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
          end
        end
        3'b001 : begin
          if(when_SuperResolutionPart1_l236) begin
            CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
          end
        end
        default : begin
        end
      endcase
    end
  end

  assign when_SuperResolutionPart1_l205 = (readStage_counterOnePixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart1_l209 = (readStage_counterTwoPixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart1_l213 = (readStage_mainTwoPixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart1_l217 = (readStage_mainOnePixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart1_l228 = (readStage_mainTwoPixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart1_l230 = (readStage_counterOnePixelStream_payload <= readStage_counterTwoPixelStream_payload);
  assign when_SuperResolutionPart1_l234 = (readStage_mainOnePixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart1_l236 = (readStage_counterTwoPixelStream_payload <= readStage_counterOnePixelStream_payload);
  assign when_SuperResolutionPart1_l241 = (readStage_counterTwoPixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart1_l246 = (readStage_counterOnePixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign readStage_controlPipe_translated_valid = readStage_controlPipe_valid;
  assign readStage_controlPipe_ready = readStage_controlPipe_translated_ready;
  assign readStage_controlPipe_translated_payload_frameStart = readStage_controlPipe_payload_frameStart;
  assign readStage_controlPipe_translated_payload_rowEnd = readStage_controlPipe_payload_rowEnd;
  assign readStage_controlPipe_translated_payload_passMode = readStage_controlPipe_payload_passMode;
  assign readStage_controlPipe_translated_payload_passValid = readStage_controlPipe_payload_passValid;
  assign readStage_controlPipe_translated_payload_onceMode = readStage_controlPipe_payload_onceMode;
  assign readStage_controlPipe_translated_payload_onceValid = readStage_controlPipe_payload_onceValid;
  assign readStage_controlPipe_translated_payload_mainCompare = CICC1851_readStage_controlPipe_translated_payload_mainCompare;
  assign readStage_controlPipe_translated_payload_counterCompare = CICC1851_readStage_controlPipe_translated_payload_counterCompare;
  assign readStage_controlPipe_translated_payload_mainDiff = readStage_controlPipe_payload_mainDiff;
  assign readStage_controlPipe_translated_payload_counterDiff = readStage_controlPipe_payload_counterDiff;
  assign readStage_controlPipe_translated_payload_twiceCompValid = readStage_controlPipe_payload_twiceCompValid;
  assign readStage_controlPipe_translated_payload_twiceMode = readStage_controlPipe_payload_twiceMode;
  assign readStage_controlPipe_translated_ready = (! readStage_controlPipe_translated_rValid);
  assign readStage_controlPipe_translated_s2mPipe_valid = (readStage_controlPipe_translated_valid || readStage_controlPipe_translated_rValid);
  assign readStage_controlPipe_translated_s2mPipe_payload_frameStart = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_frameStart : readStage_controlPipe_translated_payload_frameStart);
  assign readStage_controlPipe_translated_s2mPipe_payload_rowEnd = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_rowEnd : readStage_controlPipe_translated_payload_rowEnd);
  assign readStage_controlPipe_translated_s2mPipe_payload_passMode = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_passMode : readStage_controlPipe_translated_payload_passMode);
  assign readStage_controlPipe_translated_s2mPipe_payload_passValid = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_passValid : readStage_controlPipe_translated_payload_passValid);
  assign readStage_controlPipe_translated_s2mPipe_payload_onceMode = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_onceMode : readStage_controlPipe_translated_payload_onceMode);
  assign readStage_controlPipe_translated_s2mPipe_payload_onceValid = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_onceValid : readStage_controlPipe_translated_payload_onceValid);
  assign readStage_controlPipe_translated_s2mPipe_payload_mainCompare = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_mainCompare : readStage_controlPipe_translated_payload_mainCompare);
  assign readStage_controlPipe_translated_s2mPipe_payload_counterCompare = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_counterCompare : readStage_controlPipe_translated_payload_counterCompare);
  assign readStage_controlPipe_translated_s2mPipe_payload_mainDiff = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_mainDiff : readStage_controlPipe_translated_payload_mainDiff);
  assign readStage_controlPipe_translated_s2mPipe_payload_counterDiff = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_counterDiff : readStage_controlPipe_translated_payload_counterDiff);
  assign readStage_controlPipe_translated_s2mPipe_payload_twiceCompValid = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_twiceCompValid : readStage_controlPipe_translated_payload_twiceCompValid);
  assign readStage_controlPipe_translated_s2mPipe_payload_twiceMode = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_twiceMode : readStage_controlPipe_translated_payload_twiceMode);
  always @(*) begin
    readStage_controlPipe_translated_s2mPipe_ready = compareStage_controlPipe_ready;
    if(when_Stream_l368_15) begin
      readStage_controlPipe_translated_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_15 = (! compareStage_controlPipe_valid);
  assign compareStage_controlPipe_valid = readStage_controlPipe_translated_s2mPipe_rValid;
  assign compareStage_controlPipe_payload_frameStart = readStage_controlPipe_translated_s2mPipe_rData_frameStart;
  assign compareStage_controlPipe_payload_rowEnd = readStage_controlPipe_translated_s2mPipe_rData_rowEnd;
  assign compareStage_controlPipe_payload_passMode = readStage_controlPipe_translated_s2mPipe_rData_passMode;
  assign compareStage_controlPipe_payload_passValid = readStage_controlPipe_translated_s2mPipe_rData_passValid;
  assign compareStage_controlPipe_payload_onceMode = readStage_controlPipe_translated_s2mPipe_rData_onceMode;
  assign compareStage_controlPipe_payload_onceValid = readStage_controlPipe_translated_s2mPipe_rData_onceValid;
  assign compareStage_controlPipe_payload_mainCompare = readStage_controlPipe_translated_s2mPipe_rData_mainCompare;
  assign compareStage_controlPipe_payload_counterCompare = readStage_controlPipe_translated_s2mPipe_rData_counterCompare;
  assign compareStage_controlPipe_payload_mainDiff = readStage_controlPipe_translated_s2mPipe_rData_mainDiff;
  assign compareStage_controlPipe_payload_counterDiff = readStage_controlPipe_translated_s2mPipe_rData_counterDiff;
  assign compareStage_controlPipe_payload_twiceCompValid = readStage_controlPipe_translated_s2mPipe_rData_twiceCompValid;
  assign compareStage_controlPipe_payload_twiceMode = readStage_controlPipe_translated_s2mPipe_rData_twiceMode;
  assign compareStage_mainOnePixelStream_ready = (! compareStage_mainOnePixelStream_rValid);
  assign compareStage_mainOnePixelStream_s2mPipe_valid = (compareStage_mainOnePixelStream_valid || compareStage_mainOnePixelStream_rValid);
  assign compareStage_mainOnePixelStream_s2mPipe_payload = (compareStage_mainOnePixelStream_rValid ? compareStage_mainOnePixelStream_rData : compareStage_mainOnePixelStream_payload);
  always @(*) begin
    compareStage_mainOnePixelStream_s2mPipe_ready = diffStage_mainOnePixelStream_ready;
    if(when_Stream_l368_16) begin
      compareStage_mainOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_16 = (! diffStage_mainOnePixelStream_valid);
  assign diffStage_mainOnePixelStream_valid = compareStage_mainOnePixelStream_s2mPipe_rValid;
  assign diffStage_mainOnePixelStream_payload = compareStage_mainOnePixelStream_s2mPipe_rData;
  assign compareStage_counterOnePixelStream_ready = (! compareStage_counterOnePixelStream_rValid);
  assign compareStage_counterOnePixelStream_s2mPipe_valid = (compareStage_counterOnePixelStream_valid || compareStage_counterOnePixelStream_rValid);
  assign compareStage_counterOnePixelStream_s2mPipe_payload = (compareStage_counterOnePixelStream_rValid ? compareStage_counterOnePixelStream_rData : compareStage_counterOnePixelStream_payload);
  always @(*) begin
    compareStage_counterOnePixelStream_s2mPipe_ready = diffStage_counterOnePixelStream_ready;
    if(when_Stream_l368_17) begin
      compareStage_counterOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_17 = (! diffStage_counterOnePixelStream_valid);
  assign diffStage_counterOnePixelStream_valid = compareStage_counterOnePixelStream_s2mPipe_rValid;
  assign diffStage_counterOnePixelStream_payload = compareStage_counterOnePixelStream_s2mPipe_rData;
  assign compareStage_mainTwoPixelStream_ready = (! compareStage_mainTwoPixelStream_rValid);
  assign compareStage_mainTwoPixelStream_s2mPipe_valid = (compareStage_mainTwoPixelStream_valid || compareStage_mainTwoPixelStream_rValid);
  assign compareStage_mainTwoPixelStream_s2mPipe_payload = (compareStage_mainTwoPixelStream_rValid ? compareStage_mainTwoPixelStream_rData : compareStage_mainTwoPixelStream_payload);
  always @(*) begin
    compareStage_mainTwoPixelStream_s2mPipe_ready = diffStage_mainTwoPixelStream_ready;
    if(when_Stream_l368_18) begin
      compareStage_mainTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_18 = (! diffStage_mainTwoPixelStream_valid);
  assign diffStage_mainTwoPixelStream_valid = compareStage_mainTwoPixelStream_s2mPipe_rValid;
  assign diffStage_mainTwoPixelStream_payload = compareStage_mainTwoPixelStream_s2mPipe_rData;
  assign compareStage_counterTwoPixelStream_ready = (! compareStage_counterTwoPixelStream_rValid);
  assign compareStage_counterTwoPixelStream_s2mPipe_valid = (compareStage_counterTwoPixelStream_valid || compareStage_counterTwoPixelStream_rValid);
  assign compareStage_counterTwoPixelStream_s2mPipe_payload = (compareStage_counterTwoPixelStream_rValid ? compareStage_counterTwoPixelStream_rData : compareStage_counterTwoPixelStream_payload);
  always @(*) begin
    compareStage_counterTwoPixelStream_s2mPipe_ready = diffStage_counterTwoPixelStream_ready;
    if(when_Stream_l368_19) begin
      compareStage_counterTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_19 = (! diffStage_counterTwoPixelStream_valid);
  assign diffStage_counterTwoPixelStream_valid = compareStage_counterTwoPixelStream_s2mPipe_rValid;
  assign diffStage_counterTwoPixelStream_payload = compareStage_counterTwoPixelStream_s2mPipe_rData;
  always @(*) begin
    CICC1851_compareStage_controlPipe_translated_payload_mainDiff = compareStage_controlPipe_payload_mainDiff;
    if(compareStage_controlPipe_payload_onceValid) begin
      case(compareStage_controlPipe_payload_onceMode)
        3'b000 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_counterOnePixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterOnePixelStream_payload - compareStage_mainOnePixelStream_payload);
          end
        end
        3'b001 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterTwoPixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainTwoPixelStream_payload);
          end
        end
        3'b010 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_mainTwoPixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_mainOnePixelStream_payload);
          end
        end
        3'b011 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_mainOnePixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_mainTwoPixelStream_payload);
          end
        end
        3'b100 : begin
          CICC1851_compareStage_controlPipe_translated_payload_mainDiff = 8'h0;
        end
        3'b101 : begin
          CICC1851_compareStage_controlPipe_translated_payload_mainDiff = 8'h0;
        end
        default : begin
        end
      endcase
    end
    if(compareStage_controlPipe_payload_twiceCompValid) begin
      case(compareStage_controlPipe_payload_twiceMode)
        3'b000 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_mainTwoPixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_mainOnePixelStream_payload);
          end
        end
        3'b001 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_mainOnePixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_mainTwoPixelStream_payload);
          end
        end
        3'b010 : begin
          CICC1851_compareStage_controlPipe_translated_payload_mainDiff = 8'h0;
        end
        3'b011 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterTwoPixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainTwoPixelStream_payload);
          end
        end
        3'b100 : begin
          CICC1851_compareStage_controlPipe_translated_payload_mainDiff = 8'h0;
        end
        3'b101 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_counterOnePixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterOnePixelStream_payload - compareStage_mainOnePixelStream_payload);
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    CICC1851_compareStage_controlPipe_translated_payload_counterDiff = compareStage_controlPipe_payload_counterDiff;
    if(compareStage_controlPipe_payload_twiceCompValid) begin
      case(compareStage_controlPipe_payload_twiceMode)
        3'b000 : begin
          if(compareStage_controlPipe_payload_counterCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterTwoPixelStream_payload - compareStage_counterOnePixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterOnePixelStream_payload - compareStage_counterTwoPixelStream_payload);
          end
        end
        3'b001 : begin
          if(compareStage_controlPipe_payload_counterCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterOnePixelStream_payload - compareStage_counterTwoPixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterTwoPixelStream_payload - compareStage_counterOnePixelStream_payload);
          end
        end
        default : begin
        end
      endcase
    end
  end

  assign compareStage_controlPipe_translated_valid = compareStage_controlPipe_valid;
  assign compareStage_controlPipe_ready = compareStage_controlPipe_translated_ready;
  assign compareStage_controlPipe_translated_payload_frameStart = compareStage_controlPipe_payload_frameStart;
  assign compareStage_controlPipe_translated_payload_rowEnd = compareStage_controlPipe_payload_rowEnd;
  assign compareStage_controlPipe_translated_payload_passMode = compareStage_controlPipe_payload_passMode;
  assign compareStage_controlPipe_translated_payload_passValid = compareStage_controlPipe_payload_passValid;
  assign compareStage_controlPipe_translated_payload_onceMode = compareStage_controlPipe_payload_onceMode;
  assign compareStage_controlPipe_translated_payload_onceValid = compareStage_controlPipe_payload_onceValid;
  assign compareStage_controlPipe_translated_payload_mainCompare = compareStage_controlPipe_payload_mainCompare;
  assign compareStage_controlPipe_translated_payload_counterCompare = compareStage_controlPipe_payload_counterCompare;
  assign compareStage_controlPipe_translated_payload_mainDiff = CICC1851_compareStage_controlPipe_translated_payload_mainDiff;
  assign compareStage_controlPipe_translated_payload_counterDiff = CICC1851_compareStage_controlPipe_translated_payload_counterDiff;
  assign compareStage_controlPipe_translated_payload_twiceCompValid = compareStage_controlPipe_payload_twiceCompValid;
  assign compareStage_controlPipe_translated_payload_twiceMode = compareStage_controlPipe_payload_twiceMode;
  assign compareStage_controlPipe_translated_ready = (! compareStage_controlPipe_translated_rValid);
  assign compareStage_controlPipe_translated_s2mPipe_valid = (compareStage_controlPipe_translated_valid || compareStage_controlPipe_translated_rValid);
  assign compareStage_controlPipe_translated_s2mPipe_payload_frameStart = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_frameStart : compareStage_controlPipe_translated_payload_frameStart);
  assign compareStage_controlPipe_translated_s2mPipe_payload_rowEnd = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_rowEnd : compareStage_controlPipe_translated_payload_rowEnd);
  assign compareStage_controlPipe_translated_s2mPipe_payload_passMode = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_passMode : compareStage_controlPipe_translated_payload_passMode);
  assign compareStage_controlPipe_translated_s2mPipe_payload_passValid = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_passValid : compareStage_controlPipe_translated_payload_passValid);
  assign compareStage_controlPipe_translated_s2mPipe_payload_onceMode = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_onceMode : compareStage_controlPipe_translated_payload_onceMode);
  assign compareStage_controlPipe_translated_s2mPipe_payload_onceValid = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_onceValid : compareStage_controlPipe_translated_payload_onceValid);
  assign compareStage_controlPipe_translated_s2mPipe_payload_mainCompare = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_mainCompare : compareStage_controlPipe_translated_payload_mainCompare);
  assign compareStage_controlPipe_translated_s2mPipe_payload_counterCompare = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_counterCompare : compareStage_controlPipe_translated_payload_counterCompare);
  assign compareStage_controlPipe_translated_s2mPipe_payload_mainDiff = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_mainDiff : compareStage_controlPipe_translated_payload_mainDiff);
  assign compareStage_controlPipe_translated_s2mPipe_payload_counterDiff = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_counterDiff : compareStage_controlPipe_translated_payload_counterDiff);
  assign compareStage_controlPipe_translated_s2mPipe_payload_twiceCompValid = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_twiceCompValid : compareStage_controlPipe_translated_payload_twiceCompValid);
  assign compareStage_controlPipe_translated_s2mPipe_payload_twiceMode = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_twiceMode : compareStage_controlPipe_translated_payload_twiceMode);
  always @(*) begin
    compareStage_controlPipe_translated_s2mPipe_ready = diffStage_controlPipe_ready;
    if(when_Stream_l368_20) begin
      compareStage_controlPipe_translated_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_20 = (! diffStage_controlPipe_valid);
  assign diffStage_controlPipe_valid = compareStage_controlPipe_translated_s2mPipe_rValid;
  assign diffStage_controlPipe_payload_frameStart = compareStage_controlPipe_translated_s2mPipe_rData_frameStart;
  assign diffStage_controlPipe_payload_rowEnd = compareStage_controlPipe_translated_s2mPipe_rData_rowEnd;
  assign diffStage_controlPipe_payload_passMode = compareStage_controlPipe_translated_s2mPipe_rData_passMode;
  assign diffStage_controlPipe_payload_passValid = compareStage_controlPipe_translated_s2mPipe_rData_passValid;
  assign diffStage_controlPipe_payload_onceMode = compareStage_controlPipe_translated_s2mPipe_rData_onceMode;
  assign diffStage_controlPipe_payload_onceValid = compareStage_controlPipe_translated_s2mPipe_rData_onceValid;
  assign diffStage_controlPipe_payload_mainCompare = compareStage_controlPipe_translated_s2mPipe_rData_mainCompare;
  assign diffStage_controlPipe_payload_counterCompare = compareStage_controlPipe_translated_s2mPipe_rData_counterCompare;
  assign diffStage_controlPipe_payload_mainDiff = compareStage_controlPipe_translated_s2mPipe_rData_mainDiff;
  assign diffStage_controlPipe_payload_counterDiff = compareStage_controlPipe_translated_s2mPipe_rData_counterDiff;
  assign diffStage_controlPipe_payload_twiceCompValid = compareStage_controlPipe_translated_s2mPipe_rData_twiceCompValid;
  assign diffStage_controlPipe_payload_twiceMode = compareStage_controlPipe_translated_s2mPipe_rData_twiceMode;
  assign diffStage_mainOnePixelStream_ready = (! diffStage_mainOnePixelStream_rValid);
  assign diffStage_mainOnePixelStream_s2mPipe_valid = (diffStage_mainOnePixelStream_valid || diffStage_mainOnePixelStream_rValid);
  assign diffStage_mainOnePixelStream_s2mPipe_payload = (diffStage_mainOnePixelStream_rValid ? diffStage_mainOnePixelStream_rData : diffStage_mainOnePixelStream_payload);
  always @(*) begin
    diffStage_mainOnePixelStream_s2mPipe_ready = resultStage_mainOnePixelStream_ready;
    if(when_Stream_l368_21) begin
      diffStage_mainOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_21 = (! resultStage_mainOnePixelStream_valid);
  assign resultStage_mainOnePixelStream_valid = diffStage_mainOnePixelStream_s2mPipe_rValid;
  assign resultStage_mainOnePixelStream_payload = diffStage_mainOnePixelStream_s2mPipe_rData;
  assign diffStage_counterOnePixelStream_ready = (! diffStage_counterOnePixelStream_rValid);
  assign diffStage_counterOnePixelStream_s2mPipe_valid = (diffStage_counterOnePixelStream_valid || diffStage_counterOnePixelStream_rValid);
  assign diffStage_counterOnePixelStream_s2mPipe_payload = (diffStage_counterOnePixelStream_rValid ? diffStage_counterOnePixelStream_rData : diffStage_counterOnePixelStream_payload);
  always @(*) begin
    diffStage_counterOnePixelStream_s2mPipe_ready = resultStage_counterOnePixelStream_ready;
    if(when_Stream_l368_22) begin
      diffStage_counterOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_22 = (! resultStage_counterOnePixelStream_valid);
  assign resultStage_counterOnePixelStream_valid = diffStage_counterOnePixelStream_s2mPipe_rValid;
  assign resultStage_counterOnePixelStream_payload = diffStage_counterOnePixelStream_s2mPipe_rData;
  assign diffStage_mainTwoPixelStream_ready = (! diffStage_mainTwoPixelStream_rValid);
  assign diffStage_mainTwoPixelStream_s2mPipe_valid = (diffStage_mainTwoPixelStream_valid || diffStage_mainTwoPixelStream_rValid);
  assign diffStage_mainTwoPixelStream_s2mPipe_payload = (diffStage_mainTwoPixelStream_rValid ? diffStage_mainTwoPixelStream_rData : diffStage_mainTwoPixelStream_payload);
  always @(*) begin
    diffStage_mainTwoPixelStream_s2mPipe_ready = resultStage_mainTwoPixelStream_ready;
    if(when_Stream_l368_23) begin
      diffStage_mainTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_23 = (! resultStage_mainTwoPixelStream_valid);
  assign resultStage_mainTwoPixelStream_valid = diffStage_mainTwoPixelStream_s2mPipe_rValid;
  assign resultStage_mainTwoPixelStream_payload = diffStage_mainTwoPixelStream_s2mPipe_rData;
  assign diffStage_counterTwoPixelStream_ready = (! diffStage_counterTwoPixelStream_rValid);
  assign diffStage_counterTwoPixelStream_s2mPipe_valid = (diffStage_counterTwoPixelStream_valid || diffStage_counterTwoPixelStream_rValid);
  assign diffStage_counterTwoPixelStream_s2mPipe_payload = (diffStage_counterTwoPixelStream_rValid ? diffStage_counterTwoPixelStream_rData : diffStage_counterTwoPixelStream_payload);
  always @(*) begin
    diffStage_counterTwoPixelStream_s2mPipe_ready = resultStage_counterTwoPixelStream_ready;
    if(when_Stream_l368_24) begin
      diffStage_counterTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_24 = (! resultStage_counterTwoPixelStream_valid);
  assign resultStage_counterTwoPixelStream_valid = diffStage_counterTwoPixelStream_s2mPipe_rValid;
  assign resultStage_counterTwoPixelStream_payload = diffStage_counterTwoPixelStream_s2mPipe_rData;
  assign diffStage_controlPipe_ready = diffStage_controlPipe_fork_io_input_ready;
  assign diffStage_controlPipe_fork_io_outputs_0_ready = (! diffStage_controlPipe_fork_io_outputs_0_rValid);
  assign diffStage_controlPipe_fork_io_outputs_0_s2mPipe_valid = (diffStage_controlPipe_fork_io_outputs_0_valid || diffStage_controlPipe_fork_io_outputs_0_rValid);
  assign diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_frameStart = (diffStage_controlPipe_fork_io_outputs_0_rValid ? diffStage_controlPipe_fork_io_outputs_0_rData_frameStart : diffStage_controlPipe_fork_io_outputs_0_payload_frameStart);
  assign diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_rowEnd = (diffStage_controlPipe_fork_io_outputs_0_rValid ? diffStage_controlPipe_fork_io_outputs_0_rData_rowEnd : diffStage_controlPipe_fork_io_outputs_0_payload_rowEnd);
  assign diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_passMode = (diffStage_controlPipe_fork_io_outputs_0_rValid ? diffStage_controlPipe_fork_io_outputs_0_rData_passMode : diffStage_controlPipe_fork_io_outputs_0_payload_passMode);
  assign diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_passValid = (diffStage_controlPipe_fork_io_outputs_0_rValid ? diffStage_controlPipe_fork_io_outputs_0_rData_passValid : diffStage_controlPipe_fork_io_outputs_0_payload_passValid);
  assign diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_onceMode = (diffStage_controlPipe_fork_io_outputs_0_rValid ? diffStage_controlPipe_fork_io_outputs_0_rData_onceMode : diffStage_controlPipe_fork_io_outputs_0_payload_onceMode);
  assign diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_onceValid = (diffStage_controlPipe_fork_io_outputs_0_rValid ? diffStage_controlPipe_fork_io_outputs_0_rData_onceValid : diffStage_controlPipe_fork_io_outputs_0_payload_onceValid);
  assign diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_mainCompare = (diffStage_controlPipe_fork_io_outputs_0_rValid ? diffStage_controlPipe_fork_io_outputs_0_rData_mainCompare : diffStage_controlPipe_fork_io_outputs_0_payload_mainCompare);
  assign diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_counterCompare = (diffStage_controlPipe_fork_io_outputs_0_rValid ? diffStage_controlPipe_fork_io_outputs_0_rData_counterCompare : diffStage_controlPipe_fork_io_outputs_0_payload_counterCompare);
  assign diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_mainDiff = (diffStage_controlPipe_fork_io_outputs_0_rValid ? diffStage_controlPipe_fork_io_outputs_0_rData_mainDiff : diffStage_controlPipe_fork_io_outputs_0_payload_mainDiff);
  assign diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_counterDiff = (diffStage_controlPipe_fork_io_outputs_0_rValid ? diffStage_controlPipe_fork_io_outputs_0_rData_counterDiff : diffStage_controlPipe_fork_io_outputs_0_payload_counterDiff);
  assign diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_twiceCompValid = (diffStage_controlPipe_fork_io_outputs_0_rValid ? diffStage_controlPipe_fork_io_outputs_0_rData_twiceCompValid : diffStage_controlPipe_fork_io_outputs_0_payload_twiceCompValid);
  assign diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_twiceMode = (diffStage_controlPipe_fork_io_outputs_0_rValid ? diffStage_controlPipe_fork_io_outputs_0_rData_twiceMode : diffStage_controlPipe_fork_io_outputs_0_payload_twiceMode);
  always @(*) begin
    diffStage_controlPipe_fork_io_outputs_0_s2mPipe_ready = resultStage_controlPipe_ready;
    if(when_Stream_l368_25) begin
      diffStage_controlPipe_fork_io_outputs_0_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_25 = (! resultStage_controlPipe_valid);
  assign resultStage_controlPipe_valid = diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rValid;
  assign resultStage_controlPipe_payload_frameStart = diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_frameStart;
  assign resultStage_controlPipe_payload_rowEnd = diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_rowEnd;
  assign resultStage_controlPipe_payload_passMode = diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_passMode;
  assign resultStage_controlPipe_payload_passValid = diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_passValid;
  assign resultStage_controlPipe_payload_onceMode = diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_onceMode;
  assign resultStage_controlPipe_payload_onceValid = diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_onceValid;
  assign resultStage_controlPipe_payload_mainCompare = diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_mainCompare;
  assign resultStage_controlPipe_payload_counterCompare = diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_counterCompare;
  assign resultStage_controlPipe_payload_mainDiff = diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_mainDiff;
  assign resultStage_controlPipe_payload_counterDiff = diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_counterDiff;
  assign resultStage_controlPipe_payload_twiceCompValid = diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_twiceCompValid;
  assign resultStage_controlPipe_payload_twiceMode = diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_twiceMode;
  assign resultStage_pixelStream_valid = diffStage_controlPipe_fork_io_outputs_1_valid;
  always @(*) begin
    resultStage_pixelStream_payload = 8'h0;
    if(diffStage_controlPipe_fork_io_outputs_1_payload_passValid) begin
      if(diffStage_controlPipe_fork_io_outputs_1_payload_passMode) begin
        resultStage_pixelStream_payload = diffStage_mainTwoPixelStream_payload;
      end else begin
        resultStage_pixelStream_payload = diffStage_mainOnePixelStream_payload;
      end
    end
    if(diffStage_controlPipe_fork_io_outputs_1_payload_onceValid) begin
      case(diffStage_controlPipe_fork_io_outputs_1_payload_onceMode)
        3'b000 : begin
          if(when_SuperResolutionPart1_l339) begin
            resultStage_pixelStream_payload = diffStage_mainOnePixelStream_payload;
          end else begin
            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload[7:0];
          end
        end
        3'b001 : begin
          if(when_SuperResolutionPart1_l343) begin
            resultStage_pixelStream_payload = diffStage_mainTwoPixelStream_payload;
          end else begin
            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_2[7:0];
          end
        end
        3'b010 : begin
          if(when_SuperResolutionPart1_l347) begin
            resultStage_pixelStream_payload = diffStage_mainOnePixelStream_payload;
          end else begin
            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_4[7:0];
          end
        end
        3'b011 : begin
          if(when_SuperResolutionPart1_l351) begin
            resultStage_pixelStream_payload = diffStage_mainTwoPixelStream_payload;
          end else begin
            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_6[7:0];
          end
        end
        3'b100 : begin
          resultStage_pixelStream_payload = diffStage_mainTwoPixelStream_payload;
        end
        3'b101 : begin
          resultStage_pixelStream_payload = diffStage_mainOnePixelStream_payload;
        end
        default : begin
        end
      endcase
    end
    if(diffStage_controlPipe_fork_io_outputs_1_payload_twiceCompValid) begin
      case(diffStage_controlPipe_fork_io_outputs_1_payload_twiceMode)
        3'b000 : begin
          if(when_SuperResolutionPart1_l362) begin
            if(when_SuperResolutionPart1_l363) begin
              resultStage_pixelStream_payload = diffStage_mainOnePixelStream_payload;
            end else begin
              resultStage_pixelStream_payload = diffStage_counterTwoPixelStream_payload;
            end
          end else begin
            if(when_SuperResolutionPart1_l366) begin
              resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_8[7:0];
            end else begin
              resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_10[7:0];
            end
          end
        end
        3'b001 : begin
          if(when_SuperResolutionPart1_l371) begin
            if(when_SuperResolutionPart1_l372) begin
              resultStage_pixelStream_payload = diffStage_mainTwoPixelStream_payload;
            end else begin
              resultStage_pixelStream_payload = diffStage_counterOnePixelStream_payload;
            end
          end else begin
            if(when_SuperResolutionPart1_l375) begin
              resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_12[7:0];
            end else begin
              resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_14[7:0];
            end
          end
        end
        3'b010 : begin
          resultStage_pixelStream_payload = diffStage_mainTwoPixelStream_payload;
        end
        3'b011 : begin
          if(when_SuperResolutionPart1_l381) begin
            resultStage_pixelStream_payload = diffStage_mainTwoPixelStream_payload;
          end else begin
            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_16[7:0];
          end
        end
        3'b100 : begin
          resultStage_pixelStream_payload = diffStage_mainOnePixelStream_payload;
        end
        3'b101 : begin
          if(when_SuperResolutionPart1_l386) begin
            resultStage_pixelStream_payload = diffStage_mainOnePixelStream_payload;
          end else begin
            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_18[7:0];
          end
        end
        default : begin
        end
      endcase
    end
  end

  assign when_SuperResolutionPart1_l339 = (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart1_l343 = (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart1_l347 = (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart1_l351 = (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart1_l362 = ((inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff) && (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff));
  assign when_SuperResolutionPart1_l363 = (diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart1_l366 = (diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart1_l371 = ((inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff) && (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff));
  assign when_SuperResolutionPart1_l372 = (diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart1_l375 = (diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart1_l381 = (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart1_l386 = (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign resultStage_pixelStream_ready = (! resultStage_pixelStream_rValid);
  assign resultStage_pixelStream_s2mPipe_valid = (resultStage_pixelStream_valid || resultStage_pixelStream_rValid);
  assign resultStage_pixelStream_s2mPipe_payload = (resultStage_pixelStream_rValid ? resultStage_pixelStream_rData : resultStage_pixelStream_payload);
  always @(*) begin
    resultStage_pixelStream_s2mPipe_ready = resultStage_resultStream_ready;
    if(when_Stream_l368_26) begin
      resultStage_pixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_26 = (! resultStage_resultStream_valid);
  assign resultStage_resultStream_valid = resultStage_pixelStream_s2mPipe_rValid;
  assign resultStage_resultStream_payload = resultStage_pixelStream_s2mPipe_rData;
  assign CICC1851_resultStage_mainOnePixelStream_ready_2 = (CICC1851_resultStage_mainOnePixelStream_ready && CICC1851_resultStage_mainOnePixelStream_ready_1);
  assign CICC1851_resultStage_mainOnePixelStream_ready = (((((resultStage_resultStream_valid && resultStage_mainOnePixelStream_valid) && resultStage_counterOnePixelStream_valid) && resultStage_mainTwoPixelStream_valid) && resultStage_counterTwoPixelStream_valid) && resultStage_controlPipe_valid);
  assign resultStage_resultStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_mainOnePixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_counterOnePixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_mainTwoPixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_counterTwoPixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_controlPipe_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign when_Stream_l438 = (((! resultStage_controlPipe_payload_passValid) && (! resultStage_controlPipe_payload_onceValid)) && (! resultStage_controlPipe_payload_twiceCompValid));
  always @(*) begin
    resultsJoin_valid = CICC1851_resultStage_mainOnePixelStream_ready;
    if(when_Stream_l438) begin
      resultsJoin_valid = 1'b0;
    end
  end

  always @(*) begin
    CICC1851_resultStage_mainOnePixelStream_ready_1 = resultsJoin_ready;
    if(when_Stream_l438) begin
      CICC1851_resultStage_mainOnePixelStream_ready_1 = 1'b1;
    end
  end

  assign pixelsStream_valid = resultsJoin_valid;
  assign resultsJoin_ready = pixelsStream_ready;
  assign pixelsStream_payload_pixel = resultStage_resultStream_payload;
  assign pixelsStream_payload_frameStart = resultStage_controlPipe_payload_frameStart;
  assign pixelsStream_payload_rowEnd = resultStage_controlPipe_payload_rowEnd;
  assign pixelsStream_ready = (! pixelsStream_rValid);
  assign pixelsStream_s2mPipe_valid = (pixelsStream_valid || pixelsStream_rValid);
  assign pixelsStream_s2mPipe_payload_pixel = (pixelsStream_rValid ? pixelsStream_rData_pixel : pixelsStream_payload_pixel);
  assign pixelsStream_s2mPipe_payload_frameStart = (pixelsStream_rValid ? pixelsStream_rData_frameStart : pixelsStream_payload_frameStart);
  assign pixelsStream_s2mPipe_payload_rowEnd = (pixelsStream_rValid ? pixelsStream_rData_rowEnd : pixelsStream_payload_rowEnd);
  always @(*) begin
    pixelsStream_s2mPipe_ready = pixelsStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_27) begin
      pixelsStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_27 = (! pixelsStream_s2mPipe_m2sPipe_valid);
  assign pixelsStream_s2mPipe_m2sPipe_valid = pixelsStream_s2mPipe_rValid;
  assign pixelsStream_s2mPipe_m2sPipe_payload_pixel = pixelsStream_s2mPipe_rData_pixel;
  assign pixelsStream_s2mPipe_m2sPipe_payload_frameStart = pixelsStream_s2mPipe_rData_frameStart;
  assign pixelsStream_s2mPipe_m2sPipe_payload_rowEnd = pixelsStream_s2mPipe_rData_rowEnd;
  assign pixelsStream_s2mPipe_m2sPipe_ready = pixelsOut_ready;
  assign pixelsIn_s2mPipe_valid = (pixelsIn_valid || pixelsIn_rValid);
  assign pixelsIn_s2mPipe_payload_pixel = (pixelsIn_rValid ? pixelsIn_rData_pixel : pixelsIn_payload_pixel);
  assign pixelsIn_s2mPipe_payload_frameStart = (pixelsIn_rValid ? pixelsIn_rData_frameStart : pixelsIn_payload_frameStart);
  assign pixelsIn_s2mPipe_payload_rowEnd = (pixelsIn_rValid ? pixelsIn_rData_rowEnd : pixelsIn_payload_rowEnd);
  always @(*) begin
    pixelsIn_s2mPipe_ready = pixelsIn_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_28) begin
      pixelsIn_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_28 = (! pixelsIn_s2mPipe_m2sPipe_valid);
  assign pixelsIn_s2mPipe_m2sPipe_valid = pixelsIn_s2mPipe_rValid;
  assign pixelsIn_s2mPipe_m2sPipe_payload_pixel = pixelsIn_s2mPipe_rData_pixel;
  assign pixelsIn_s2mPipe_m2sPipe_payload_frameStart = pixelsIn_s2mPipe_rData_frameStart;
  assign pixelsIn_s2mPipe_m2sPipe_payload_rowEnd = pixelsIn_s2mPipe_rData_rowEnd;
  assign passPixels_valid = (pixelsIn_s2mPipe_m2sPipe_valid && bufferEnable);
  assign pixelsIn_s2mPipe_m2sPipe_ready = (passPixels_ready && bufferEnable);
  assign passPixels_payload_pixel = pixelsIn_s2mPipe_m2sPipe_payload_pixel;
  assign passPixels_payload_frameStart = pixelsIn_s2mPipe_m2sPipe_payload_frameStart;
  assign passPixels_payload_rowEnd = pixelsIn_s2mPipe_m2sPipe_payload_rowEnd;
  assign passPixels_ready = 1'b1;
  assign passPixels_fire = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart1_l421 = ((bufferWAddr_value == CICC1851_when_SuperResolutionPart1_l421) && passPixels_fire);
  assign passPixels_fire_1 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart1_l422 = (((bufferRowCount_value == CICC1851_when_SuperResolutionPart1_l422) && bufferReachRowEnd) && passPixels_fire_1);
  assign passPixels_fire_2 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart1_l425 = (passPixels_payload_rowEnd && passPixels_fire_2);
  assign passPixels_fire_3 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart1_l438 = (passPixels_payload_rowEnd && passPixels_fire_3);
  assign passPixels_fire_4 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart1_l439 = (((bufferRowCount_value != 10'h0) && passPixels_payload_rowEnd) && passPixels_fire_4);
  assign when_SuperResolutionPart1_l442 = (bufferReachFinalRow && bufferReachRowEnd);
  assign controlStream_fire = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l447 = (((CICC1851_when_SuperResolutionPart1_l447 == 11'h001) && controlStream_payload_rowEnd) && controlStream_fire);
  assign when_SuperResolutionPart1_l449 = 1'b1;
  assign passPixels_fire_5 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart1_l453 = (passPixels_payload_frameStart && passPixels_fire_5);
  assign passPixels_fire_6 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_7 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_8 = (passPixels_valid && passPixels_ready);
  assign controlStateMachine_wantExit = 1'b0;
  always @(*) begin
    controlStateMachine_wantStart = 1'b0;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_3_HOLD : begin
      end
      controlStateMachine_enumDef_3_PASS : begin
      end
      controlStateMachine_enumDef_3_ONCE : begin
      end
      controlStateMachine_enumDef_3_TWICE : begin
      end
      default : begin
        controlStateMachine_wantStart = 1'b1;
      end
    endcase
  end

  assign controlStateMachine_wantKill = 1'b0;
  always @(*) begin
    controlStateMachine_stateNext = controlStateMachine_stateReg;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_3_HOLD : begin
        if(when_SuperResolutionPart1_l482) begin
          if(passPixels_fire_9) begin
            if(when_SuperResolutionPart1_l484) begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_3_PASS;
            end else begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_3_ONCE;
            end
          end
        end else begin
          if(passPixels_fire_10) begin
            if(when_SuperResolutionPart1_l489) begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_3_ONCE;
            end else begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_3_TWICE;
            end
          end
        end
      end
      controlStateMachine_enumDef_3_PASS : begin
        if(controlStream_fire_1) begin
          if(when_SuperResolutionPart1_l498) begin
            controlStateMachine_stateNext = controlStateMachine_enumDef_3_ONCE;
          end else begin
            if(when_SuperResolutionPart1_l500) begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_3_HOLD;
            end else begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_3_ONCE;
            end
          end
        end
      end
      controlStateMachine_enumDef_3_ONCE : begin
        if(when_SuperResolutionPart1_l537) begin
          if(controlStream_fire_7) begin
            if(outReachRowEnd) begin
              if(bufferReuse) begin
                controlStateMachine_stateNext = controlStateMachine_enumDef_3_ONCE;
              end else begin
                if(when_SuperResolutionPart1_l542) begin
                  controlStateMachine_stateNext = controlStateMachine_enumDef_3_HOLD;
                end else begin
                  controlStateMachine_stateNext = controlStateMachine_enumDef_3_ONCE;
                end
              end
            end else begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_3_PASS;
            end
          end
        end else begin
          if(controlStream_fire_8) begin
            if(bufferReuse) begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_3_TWICE;
            end else begin
              if(when_SuperResolutionPart1_l563) begin
                controlStateMachine_stateNext = controlStateMachine_enumDef_3_HOLD;
              end else begin
                controlStateMachine_stateNext = controlStateMachine_enumDef_3_TWICE;
              end
            end
          end
        end
      end
      controlStateMachine_enumDef_3_TWICE : begin
        if(controlStream_fire_13) begin
          if(outReachRowEnd) begin
            if(bufferReuse) begin
              if(outReachFinalRow) begin
                controlStateMachine_stateNext = controlStateMachine_enumDef_3_HOLD;
              end else begin
                controlStateMachine_stateNext = controlStateMachine_enumDef_3_PASS;
              end
            end else begin
              if(when_SuperResolutionPart1_l612) begin
                controlStateMachine_stateNext = controlStateMachine_enumDef_3_HOLD;
              end else begin
                controlStateMachine_stateNext = controlStateMachine_enumDef_3_PASS;
              end
            end
          end else begin
            controlStateMachine_stateNext = controlStateMachine_enumDef_3_ONCE;
          end
        end
      end
      default : begin
      end
    endcase
    if(controlStateMachine_wantStart) begin
      controlStateMachine_stateNext = controlStateMachine_enumDef_3_HOLD;
    end
    if(controlStateMachine_wantKill) begin
      controlStateMachine_stateNext = controlStateMachine_enumDef_3_BOOT;
    end
  end

  assign when_SuperResolutionPart1_l482 = (CICC1851_when_SuperResolutionPart1_l482 == 11'h0);
  assign passPixels_fire_9 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart1_l484 = (CICC1851_when_SuperResolutionPart1_l484 == 11'h0);
  assign passPixels_fire_10 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart1_l489 = (CICC1851_when_SuperResolutionPart1_l489 == 11'h0);
  assign controlStream_fire_1 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l498 = ((CICC1851_when_SuperResolutionPart1_l498 < CICC1851_when_SuperResolutionPart1_l498_1) || bufferReuse);
  assign passPixels_fire_11 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart1_l500 = ((CICC1851_when_SuperResolutionPart1_l500 == CICC1851_when_SuperResolutionPart1_l500_1) && (! passPixels_fire_11));
  assign controlStream_fire_2 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l507 = (frameStart && controlStream_fire_2);
  assign controlStream_fire_3 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l510 = (controlStream_fire_3 && (CICC1851_when_SuperResolutionPart1_l510 == CICC1851_when_SuperResolutionPart1_l510_1));
  assign controlStream_fire_4 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l511 = ((outReachRowEnd && (CICC1851_when_SuperResolutionPart1_l511 == CICC1851_when_SuperResolutionPart1_l511_1)) && controlStream_fire_4);
  assign controlStream_fire_5 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l513 = (controlStream_fire_5 && outReachRowEnd);
  assign controlStream_fire_6 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l537 = (CICC1851_when_SuperResolutionPart1_l537 == 11'h0);
  assign controlStream_fire_7 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l542 = ((bufferWAddr_value == 10'h0) && (CICC1851_when_SuperResolutionPart1_l542 == CICC1851_when_SuperResolutionPart1_l542_2));
  assign controlStream_fire_8 = (controlStream_valid && controlStream_ready);
  assign passPixels_fire_12 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart1_l563 = ((CICC1851_when_SuperResolutionPart1_l563 == CICC1851_when_SuperResolutionPart1_l563_1) && (! passPixels_fire_12));
  assign controlStream_fire_9 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l578 = (controlStream_fire_9 && (CICC1851_when_SuperResolutionPart1_l578 == CICC1851_when_SuperResolutionPart1_l578_1));
  assign controlStream_fire_10 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l579 = ((outReachRowEnd && (CICC1851_when_SuperResolutionPart1_l579 == CICC1851_when_SuperResolutionPart1_l579_1)) && controlStream_fire_10);
  assign controlStream_fire_11 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l581 = (controlStream_fire_11 && outReachRowEnd);
  assign controlStream_fire_12 = (controlStream_valid && controlStream_ready);
  assign controlStream_fire_13 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l612 = (bufferWAddr_value == 10'h0);
  assign controlStream_fire_14 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l664 = (controlStream_fire_14 && (CICC1851_when_SuperResolutionPart1_l664 == CICC1851_when_SuperResolutionPart1_l664_1));
  assign controlStream_fire_15 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l665 = ((outReachRowEnd && (CICC1851_when_SuperResolutionPart1_l665 == CICC1851_when_SuperResolutionPart1_l665_1)) && controlStream_fire_15);
  assign controlStream_fire_16 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l667 = (controlStream_fire_16 && outReachRowEnd);
  assign controlStream_fire_17 = (controlStream_valid && controlStream_ready);
  always @(posedge clk or negedge resetn) begin
    if(!resetn) begin
      inpDone <= 1'b0;
      readDone <= 1'b0;
      startRead <= 1'b0;
      slaveStart <= 1'b0;
      frameStart <= 1'b0;
      inpThreshold <= 8'h80;
      bmpWidth <= 10'h3c0;
      bmpHeight <= 10'h21c;
      holdBuffer <= 1'b0;
      writeDone <= 1'b0;
      bufferRowCount_value <= 10'h0;
      bufferEnable <= 1'b0;
      bufferSwitch <= 1'b0;
      nextRowBuffer <= 1'b1;
      bufferReuse <= 1'b0;
      bufferWAddr_value <= 10'h0;
      outPixelAddr_value <= 11'h0;
      outRowCount_value <= 11'h0;
      outReachRowEnd <= 1'b0;
      outReachFinalRow <= 1'b0;
      bufferReachRowEnd <= 1'b0;
      bufferReachFinalRow <= 1'b0;
      mainAddrOneStream_rValid <= 1'b0;
      mainAddrOneStream_s2mPipe_rValid <= 1'b0;
      CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_mainOnePixelStream_valid <= 1'b0;
      counterAddrOneStream_rValid <= 1'b0;
      counterAddrOneStream_s2mPipe_rValid <= 1'b0;
      CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_counterOnePixelStream_valid <= 1'b0;
      mainAddrTwoStream_rValid <= 1'b0;
      mainAddrTwoStream_s2mPipe_rValid <= 1'b0;
      CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_mainTwoPixelStream_valid <= 1'b0;
      counterAddrTwoStream_rValid <= 1'b0;
      counterAddrTwoStream_s2mPipe_rValid <= 1'b0;
      CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_counterTwoPixelStream_valid <= 1'b0;
      controlStream_rValid <= 1'b0;
      controlStream_s2mPipe_rValid <= 1'b0;
      controlStream_s2mPipe_m2sPipe_rValid <= 1'b0;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rValid <= 1'b0;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rValid <= 1'b0;
      readStage_mainOnePixelStream_rValid <= 1'b0;
      readStage_mainOnePixelStream_s2mPipe_rValid <= 1'b0;
      readStage_counterOnePixelStream_rValid <= 1'b0;
      readStage_counterOnePixelStream_s2mPipe_rValid <= 1'b0;
      readStage_mainTwoPixelStream_rValid <= 1'b0;
      readStage_mainTwoPixelStream_s2mPipe_rValid <= 1'b0;
      readStage_counterTwoPixelStream_rValid <= 1'b0;
      readStage_counterTwoPixelStream_s2mPipe_rValid <= 1'b0;
      readStage_controlPipe_translated_rValid <= 1'b0;
      readStage_controlPipe_translated_s2mPipe_rValid <= 1'b0;
      compareStage_mainOnePixelStream_rValid <= 1'b0;
      compareStage_mainOnePixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_counterOnePixelStream_rValid <= 1'b0;
      compareStage_counterOnePixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_mainTwoPixelStream_rValid <= 1'b0;
      compareStage_mainTwoPixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_counterTwoPixelStream_rValid <= 1'b0;
      compareStage_counterTwoPixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_controlPipe_translated_rValid <= 1'b0;
      compareStage_controlPipe_translated_s2mPipe_rValid <= 1'b0;
      diffStage_mainOnePixelStream_rValid <= 1'b0;
      diffStage_mainOnePixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_counterOnePixelStream_rValid <= 1'b0;
      diffStage_counterOnePixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_mainTwoPixelStream_rValid <= 1'b0;
      diffStage_mainTwoPixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_counterTwoPixelStream_rValid <= 1'b0;
      diffStage_counterTwoPixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_controlPipe_fork_io_outputs_0_rValid <= 1'b0;
      diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rValid <= 1'b0;
      resultStage_pixelStream_rValid <= 1'b0;
      resultStage_pixelStream_s2mPipe_rValid <= 1'b0;
      pixelsStream_rValid <= 1'b0;
      pixelsStream_s2mPipe_rValid <= 1'b0;
      pixelsIn_rValid <= 1'b0;
      pixelsIn_s2mPipe_rValid <= 1'b0;
      controlStateMachine_stateReg <= controlStateMachine_enumDef_3_BOOT;
    end else begin
      if(when_SuperResolutionPart1_l79) begin
        inpDone <= 1'b1;
      end
      if(when_SuperResolutionPart1_l79_1) begin
        inpDone <= 1'b0;
      end
      if(when_SuperResolutionPart1_l82) begin
        readDone <= 1'b0;
      end
      if(when_SuperResolutionPart1_l85) begin
        startRead <= 1'b1;
      end
      if(when_SuperResolutionPart1_l85_1) begin
        startRead <= 1'b0;
      end
      if(when_SuperResolutionPart1_l88) begin
        slaveStart <= 1'b1;
      end
      if(when_SuperResolutionPart1_l88_1) begin
        slaveStart <= 1'b0;
      end
      inpThreshold <= thresholdIn;
      bmpWidth <= widthIn;
      bmpHeight <= heightIn;
      if(when_SuperResolutionPart1_l103) begin
        holdBuffer <= 1'b0;
      end
      if(when_SuperResolutionPart1_l106) begin
        writeDone <= 1'b0;
      end
      bufferRowCount_value <= bufferRowCount_valueNext;
      if(when_SuperResolutionPart1_l112) begin
        bufferEnable <= 1'b1;
      end
      if(when_SuperResolutionPart1_l112_1) begin
        bufferEnable <= 1'b0;
      end
      if(when_SuperResolutionPart1_l115) begin
        bufferSwitch <= 1'b0;
      end
      if(when_SuperResolutionPart1_l118) begin
        nextRowBuffer <= 1'b1;
      end
      if(inpDone) begin
        bufferReuse <= 1'b0;
      end
      bufferWAddr_value <= bufferWAddr_valueNext;
      outPixelAddr_value <= outPixelAddr_valueNext;
      outRowCount_value <= outRowCount_valueNext;
      if(mainAddrOneStream_valid) begin
        mainAddrOneStream_rValid <= 1'b1;
      end
      if(mainAddrOneStream_s2mPipe_ready) begin
        mainAddrOneStream_rValid <= 1'b0;
      end
      if(mainAddrOneStream_s2mPipe_ready) begin
        mainAddrOneStream_s2mPipe_rValid <= mainAddrOneStream_s2mPipe_valid;
      end
      if(CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(mainAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_2 <= mainAddrOneStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_1) begin
        CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_1) begin
        CICC1851_readStage_mainOnePixelStream_valid <= (CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready || CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_3);
      end
      if(counterAddrOneStream_valid) begin
        counterAddrOneStream_rValid <= 1'b1;
      end
      if(counterAddrOneStream_s2mPipe_ready) begin
        counterAddrOneStream_rValid <= 1'b0;
      end
      if(counterAddrOneStream_s2mPipe_ready) begin
        counterAddrOneStream_s2mPipe_rValid <= counterAddrOneStream_s2mPipe_valid;
      end
      if(CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(counterAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_2 <= counterAddrOneStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_2) begin
        CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_2) begin
        CICC1851_readStage_counterOnePixelStream_valid <= (CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready || CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_3);
      end
      if(mainAddrTwoStream_valid) begin
        mainAddrTwoStream_rValid <= 1'b1;
      end
      if(mainAddrTwoStream_s2mPipe_ready) begin
        mainAddrTwoStream_rValid <= 1'b0;
      end
      if(mainAddrTwoStream_s2mPipe_ready) begin
        mainAddrTwoStream_s2mPipe_rValid <= mainAddrTwoStream_s2mPipe_valid;
      end
      if(CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(mainAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= mainAddrTwoStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_3) begin
        CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_3) begin
        CICC1851_readStage_mainTwoPixelStream_valid <= (CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready || CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_3);
      end
      if(counterAddrTwoStream_valid) begin
        counterAddrTwoStream_rValid <= 1'b1;
      end
      if(counterAddrTwoStream_s2mPipe_ready) begin
        counterAddrTwoStream_rValid <= 1'b0;
      end
      if(counterAddrTwoStream_s2mPipe_ready) begin
        counterAddrTwoStream_s2mPipe_rValid <= counterAddrTwoStream_s2mPipe_valid;
      end
      if(CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(counterAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= counterAddrTwoStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_4) begin
        CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_4) begin
        CICC1851_readStage_counterTwoPixelStream_valid <= (CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready || CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_3);
      end
      if(controlStream_valid) begin
        controlStream_rValid <= 1'b1;
      end
      if(controlStream_s2mPipe_ready) begin
        controlStream_rValid <= 1'b0;
      end
      if(controlStream_s2mPipe_ready) begin
        controlStream_s2mPipe_rValid <= controlStream_s2mPipe_valid;
      end
      if(controlStream_s2mPipe_m2sPipe_ready) begin
        controlStream_s2mPipe_m2sPipe_rValid <= controlStream_s2mPipe_m2sPipe_valid;
      end
      if(controlStream_s2mPipe_m2sPipe_m2sPipe_valid) begin
        controlStream_s2mPipe_m2sPipe_m2sPipe_rValid <= 1'b1;
      end
      if(controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready) begin
        controlStream_s2mPipe_m2sPipe_m2sPipe_rValid <= 1'b0;
      end
      if(controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready) begin
        controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_valid;
      end
      if(readStage_mainOnePixelStream_valid) begin
        readStage_mainOnePixelStream_rValid <= 1'b1;
      end
      if(readStage_mainOnePixelStream_s2mPipe_ready) begin
        readStage_mainOnePixelStream_rValid <= 1'b0;
      end
      if(readStage_mainOnePixelStream_s2mPipe_ready) begin
        readStage_mainOnePixelStream_s2mPipe_rValid <= readStage_mainOnePixelStream_s2mPipe_valid;
      end
      if(readStage_counterOnePixelStream_valid) begin
        readStage_counterOnePixelStream_rValid <= 1'b1;
      end
      if(readStage_counterOnePixelStream_s2mPipe_ready) begin
        readStage_counterOnePixelStream_rValid <= 1'b0;
      end
      if(readStage_counterOnePixelStream_s2mPipe_ready) begin
        readStage_counterOnePixelStream_s2mPipe_rValid <= readStage_counterOnePixelStream_s2mPipe_valid;
      end
      if(readStage_mainTwoPixelStream_valid) begin
        readStage_mainTwoPixelStream_rValid <= 1'b1;
      end
      if(readStage_mainTwoPixelStream_s2mPipe_ready) begin
        readStage_mainTwoPixelStream_rValid <= 1'b0;
      end
      if(readStage_mainTwoPixelStream_s2mPipe_ready) begin
        readStage_mainTwoPixelStream_s2mPipe_rValid <= readStage_mainTwoPixelStream_s2mPipe_valid;
      end
      if(readStage_counterTwoPixelStream_valid) begin
        readStage_counterTwoPixelStream_rValid <= 1'b1;
      end
      if(readStage_counterTwoPixelStream_s2mPipe_ready) begin
        readStage_counterTwoPixelStream_rValid <= 1'b0;
      end
      if(readStage_counterTwoPixelStream_s2mPipe_ready) begin
        readStage_counterTwoPixelStream_s2mPipe_rValid <= readStage_counterTwoPixelStream_s2mPipe_valid;
      end
      if(readStage_controlPipe_translated_valid) begin
        readStage_controlPipe_translated_rValid <= 1'b1;
      end
      if(readStage_controlPipe_translated_s2mPipe_ready) begin
        readStage_controlPipe_translated_rValid <= 1'b0;
      end
      if(readStage_controlPipe_translated_s2mPipe_ready) begin
        readStage_controlPipe_translated_s2mPipe_rValid <= readStage_controlPipe_translated_s2mPipe_valid;
      end
      if(compareStage_mainOnePixelStream_valid) begin
        compareStage_mainOnePixelStream_rValid <= 1'b1;
      end
      if(compareStage_mainOnePixelStream_s2mPipe_ready) begin
        compareStage_mainOnePixelStream_rValid <= 1'b0;
      end
      if(compareStage_mainOnePixelStream_s2mPipe_ready) begin
        compareStage_mainOnePixelStream_s2mPipe_rValid <= compareStage_mainOnePixelStream_s2mPipe_valid;
      end
      if(compareStage_counterOnePixelStream_valid) begin
        compareStage_counterOnePixelStream_rValid <= 1'b1;
      end
      if(compareStage_counterOnePixelStream_s2mPipe_ready) begin
        compareStage_counterOnePixelStream_rValid <= 1'b0;
      end
      if(compareStage_counterOnePixelStream_s2mPipe_ready) begin
        compareStage_counterOnePixelStream_s2mPipe_rValid <= compareStage_counterOnePixelStream_s2mPipe_valid;
      end
      if(compareStage_mainTwoPixelStream_valid) begin
        compareStage_mainTwoPixelStream_rValid <= 1'b1;
      end
      if(compareStage_mainTwoPixelStream_s2mPipe_ready) begin
        compareStage_mainTwoPixelStream_rValid <= 1'b0;
      end
      if(compareStage_mainTwoPixelStream_s2mPipe_ready) begin
        compareStage_mainTwoPixelStream_s2mPipe_rValid <= compareStage_mainTwoPixelStream_s2mPipe_valid;
      end
      if(compareStage_counterTwoPixelStream_valid) begin
        compareStage_counterTwoPixelStream_rValid <= 1'b1;
      end
      if(compareStage_counterTwoPixelStream_s2mPipe_ready) begin
        compareStage_counterTwoPixelStream_rValid <= 1'b0;
      end
      if(compareStage_counterTwoPixelStream_s2mPipe_ready) begin
        compareStage_counterTwoPixelStream_s2mPipe_rValid <= compareStage_counterTwoPixelStream_s2mPipe_valid;
      end
      if(compareStage_controlPipe_translated_valid) begin
        compareStage_controlPipe_translated_rValid <= 1'b1;
      end
      if(compareStage_controlPipe_translated_s2mPipe_ready) begin
        compareStage_controlPipe_translated_rValid <= 1'b0;
      end
      if(compareStage_controlPipe_translated_s2mPipe_ready) begin
        compareStage_controlPipe_translated_s2mPipe_rValid <= compareStage_controlPipe_translated_s2mPipe_valid;
      end
      if(diffStage_mainOnePixelStream_valid) begin
        diffStage_mainOnePixelStream_rValid <= 1'b1;
      end
      if(diffStage_mainOnePixelStream_s2mPipe_ready) begin
        diffStage_mainOnePixelStream_rValid <= 1'b0;
      end
      if(diffStage_mainOnePixelStream_s2mPipe_ready) begin
        diffStage_mainOnePixelStream_s2mPipe_rValid <= diffStage_mainOnePixelStream_s2mPipe_valid;
      end
      if(diffStage_counterOnePixelStream_valid) begin
        diffStage_counterOnePixelStream_rValid <= 1'b1;
      end
      if(diffStage_counterOnePixelStream_s2mPipe_ready) begin
        diffStage_counterOnePixelStream_rValid <= 1'b0;
      end
      if(diffStage_counterOnePixelStream_s2mPipe_ready) begin
        diffStage_counterOnePixelStream_s2mPipe_rValid <= diffStage_counterOnePixelStream_s2mPipe_valid;
      end
      if(diffStage_mainTwoPixelStream_valid) begin
        diffStage_mainTwoPixelStream_rValid <= 1'b1;
      end
      if(diffStage_mainTwoPixelStream_s2mPipe_ready) begin
        diffStage_mainTwoPixelStream_rValid <= 1'b0;
      end
      if(diffStage_mainTwoPixelStream_s2mPipe_ready) begin
        diffStage_mainTwoPixelStream_s2mPipe_rValid <= diffStage_mainTwoPixelStream_s2mPipe_valid;
      end
      if(diffStage_counterTwoPixelStream_valid) begin
        diffStage_counterTwoPixelStream_rValid <= 1'b1;
      end
      if(diffStage_counterTwoPixelStream_s2mPipe_ready) begin
        diffStage_counterTwoPixelStream_rValid <= 1'b0;
      end
      if(diffStage_counterTwoPixelStream_s2mPipe_ready) begin
        diffStage_counterTwoPixelStream_s2mPipe_rValid <= diffStage_counterTwoPixelStream_s2mPipe_valid;
      end
      if(diffStage_controlPipe_fork_io_outputs_0_valid) begin
        diffStage_controlPipe_fork_io_outputs_0_rValid <= 1'b1;
      end
      if(diffStage_controlPipe_fork_io_outputs_0_s2mPipe_ready) begin
        diffStage_controlPipe_fork_io_outputs_0_rValid <= 1'b0;
      end
      if(diffStage_controlPipe_fork_io_outputs_0_s2mPipe_ready) begin
        diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rValid <= diffStage_controlPipe_fork_io_outputs_0_s2mPipe_valid;
      end
      if(resultStage_pixelStream_valid) begin
        resultStage_pixelStream_rValid <= 1'b1;
      end
      if(resultStage_pixelStream_s2mPipe_ready) begin
        resultStage_pixelStream_rValid <= 1'b0;
      end
      if(resultStage_pixelStream_s2mPipe_ready) begin
        resultStage_pixelStream_s2mPipe_rValid <= resultStage_pixelStream_s2mPipe_valid;
      end
      if(pixelsStream_valid) begin
        pixelsStream_rValid <= 1'b1;
      end
      if(pixelsStream_s2mPipe_ready) begin
        pixelsStream_rValid <= 1'b0;
      end
      if(pixelsStream_s2mPipe_ready) begin
        pixelsStream_s2mPipe_rValid <= pixelsStream_s2mPipe_valid;
      end
      if(pixelsIn_valid) begin
        pixelsIn_rValid <= 1'b1;
      end
      if(pixelsIn_s2mPipe_ready) begin
        pixelsIn_rValid <= 1'b0;
      end
      if(pixelsIn_s2mPipe_ready) begin
        pixelsIn_s2mPipe_rValid <= pixelsIn_s2mPipe_valid;
      end
      if(when_SuperResolutionPart1_l421) begin
        bufferReachRowEnd <= 1'b1;
      end
      if(when_SuperResolutionPart1_l422) begin
        bufferReachFinalRow <= 1'b1;
      end
      if(when_SuperResolutionPart1_l425) begin
        if(bufferReachFinalRow) begin
          bufferReuse <= 1'b1;
          bufferReachRowEnd <= 1'b0;
          bufferReachFinalRow <= 1'b0;
        end else begin
          bufferReachRowEnd <= 1'b0;
        end
      end
      if(when_SuperResolutionPart1_l438) begin
        bufferSwitch <= (! bufferSwitch);
      end
      if(when_SuperResolutionPart1_l439) begin
        holdBuffer <= 1'b1;
        bufferEnable <= 1'b0;
        if(when_SuperResolutionPart1_l442) begin
          writeDone <= 1'b1;
          bufferEnable <= 1'b0;
        end
      end
      if(when_SuperResolutionPart1_l447) begin
        holdBuffer <= 1'b0;
        if(when_SuperResolutionPart1_l449) begin
          nextRowBuffer <= (! nextRowBuffer);
        end
      end
      if(when_SuperResolutionPart1_l453) begin
        frameStart <= 1'b1;
      end
      if(inpDone) begin
        inpDone <= 1'b0;
      end
      controlStateMachine_stateReg <= controlStateMachine_stateNext;
      case(controlStateMachine_stateReg)
        controlStateMachine_enumDef_3_HOLD : begin
        end
        controlStateMachine_enumDef_3_PASS : begin
          if(when_SuperResolutionPart1_l507) begin
            frameStart <= 1'b0;
          end
          if(when_SuperResolutionPart1_l510) begin
            outReachRowEnd <= 1'b1;
          end
          if(when_SuperResolutionPart1_l511) begin
            outReachFinalRow <= 1'b1;
          end
          if(when_SuperResolutionPart1_l513) begin
            if(outReachFinalRow) begin
              startRead <= 1'b0;
              readDone <= 1'b1;
              outReachRowEnd <= 1'b0;
              outReachFinalRow <= 1'b0;
            end else begin
              outReachRowEnd <= 1'b0;
            end
          end
          if(controlStream_fire_6) begin
            if(outReachRowEnd) begin
              outReachRowEnd <= 1'b0;
            end
          end
        end
        controlStateMachine_enumDef_3_ONCE : begin
          if(when_SuperResolutionPart1_l578) begin
            outReachRowEnd <= 1'b1;
          end
          if(when_SuperResolutionPart1_l579) begin
            outReachFinalRow <= 1'b1;
          end
          if(when_SuperResolutionPart1_l581) begin
            if(outReachFinalRow) begin
              startRead <= 1'b0;
              readDone <= 1'b1;
              outReachRowEnd <= 1'b0;
              outReachFinalRow <= 1'b0;
            end else begin
              outReachRowEnd <= 1'b0;
            end
          end
          if(controlStream_fire_12) begin
            if(outReachRowEnd) begin
              outReachRowEnd <= 1'b0;
            end
          end
        end
        controlStateMachine_enumDef_3_TWICE : begin
          if(when_SuperResolutionPart1_l664) begin
            outReachRowEnd <= 1'b1;
          end
          if(when_SuperResolutionPart1_l665) begin
            outReachFinalRow <= 1'b1;
          end
          if(when_SuperResolutionPart1_l667) begin
            if(outReachFinalRow) begin
              startRead <= 1'b0;
              readDone <= 1'b1;
              outReachRowEnd <= 1'b0;
              outReachFinalRow <= 1'b0;
            end else begin
              outReachRowEnd <= 1'b0;
            end
          end
          if(controlStream_fire_17) begin
            if(outReachRowEnd) begin
              outReachRowEnd <= 1'b0;
            end
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(posedge clk) begin
    startIn_regNext <= startIn;
    if(mainAddrOneStream_ready) begin
      mainAddrOneStream_rData <= mainAddrOneStream_payload;
    end
    if(mainAddrOneStream_s2mPipe_ready) begin
      mainAddrOneStream_s2mPipe_rData <= mainAddrOneStream_s2mPipe_payload;
    end
    if(CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_mainOnePixelStream_payload_1 <= CICC1851_readStage_mainOnePixelStream_payload;
    end
    if(CICC1851_1) begin
      CICC1851_readStage_mainOnePixelStream_payload_2 <= (CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_mainOnePixelStream_payload_1 : CICC1851_readStage_mainOnePixelStream_payload);
    end
    if(counterAddrOneStream_ready) begin
      counterAddrOneStream_rData <= counterAddrOneStream_payload;
    end
    if(counterAddrOneStream_s2mPipe_ready) begin
      counterAddrOneStream_s2mPipe_rData <= counterAddrOneStream_s2mPipe_payload;
    end
    if(CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_counterOnePixelStream_payload_1 <= CICC1851_readStage_counterOnePixelStream_payload;
    end
    if(CICC1851_2) begin
      CICC1851_readStage_counterOnePixelStream_payload_2 <= (CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_counterOnePixelStream_payload_1 : CICC1851_readStage_counterOnePixelStream_payload);
    end
    if(mainAddrTwoStream_ready) begin
      mainAddrTwoStream_rData <= mainAddrTwoStream_payload;
    end
    if(mainAddrTwoStream_s2mPipe_ready) begin
      mainAddrTwoStream_s2mPipe_rData <= mainAddrTwoStream_s2mPipe_payload;
    end
    if(CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_mainTwoPixelStream_payload_1 <= CICC1851_readStage_mainTwoPixelStream_payload;
    end
    if(CICC1851_3) begin
      CICC1851_readStage_mainTwoPixelStream_payload_2 <= (CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_mainTwoPixelStream_payload_1 : CICC1851_readStage_mainTwoPixelStream_payload);
    end
    if(counterAddrTwoStream_ready) begin
      counterAddrTwoStream_rData <= counterAddrTwoStream_payload;
    end
    if(counterAddrTwoStream_s2mPipe_ready) begin
      counterAddrTwoStream_s2mPipe_rData <= counterAddrTwoStream_s2mPipe_payload;
    end
    if(CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_counterTwoPixelStream_payload_1 <= CICC1851_readStage_counterTwoPixelStream_payload;
    end
    if(CICC1851_4) begin
      CICC1851_readStage_counterTwoPixelStream_payload_2 <= (CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_counterTwoPixelStream_payload_1 : CICC1851_readStage_counterTwoPixelStream_payload);
    end
    if(controlStream_ready) begin
      controlStream_rData_frameStart <= controlStream_payload_frameStart;
      controlStream_rData_rowEnd <= controlStream_payload_rowEnd;
      controlStream_rData_passMode <= controlStream_payload_passMode;
      controlStream_rData_passValid <= controlStream_payload_passValid;
      controlStream_rData_onceMode <= controlStream_payload_onceMode;
      controlStream_rData_onceValid <= controlStream_payload_onceValid;
      controlStream_rData_mainCompare <= controlStream_payload_mainCompare;
      controlStream_rData_counterCompare <= controlStream_payload_counterCompare;
      controlStream_rData_mainDiff <= controlStream_payload_mainDiff;
      controlStream_rData_counterDiff <= controlStream_payload_counterDiff;
      controlStream_rData_twiceCompValid <= controlStream_payload_twiceCompValid;
      controlStream_rData_twiceMode <= controlStream_payload_twiceMode;
    end
    if(controlStream_s2mPipe_ready) begin
      controlStream_s2mPipe_rData_frameStart <= controlStream_s2mPipe_payload_frameStart;
      controlStream_s2mPipe_rData_rowEnd <= controlStream_s2mPipe_payload_rowEnd;
      controlStream_s2mPipe_rData_passMode <= controlStream_s2mPipe_payload_passMode;
      controlStream_s2mPipe_rData_passValid <= controlStream_s2mPipe_payload_passValid;
      controlStream_s2mPipe_rData_onceMode <= controlStream_s2mPipe_payload_onceMode;
      controlStream_s2mPipe_rData_onceValid <= controlStream_s2mPipe_payload_onceValid;
      controlStream_s2mPipe_rData_mainCompare <= controlStream_s2mPipe_payload_mainCompare;
      controlStream_s2mPipe_rData_counterCompare <= controlStream_s2mPipe_payload_counterCompare;
      controlStream_s2mPipe_rData_mainDiff <= controlStream_s2mPipe_payload_mainDiff;
      controlStream_s2mPipe_rData_counterDiff <= controlStream_s2mPipe_payload_counterDiff;
      controlStream_s2mPipe_rData_twiceCompValid <= controlStream_s2mPipe_payload_twiceCompValid;
      controlStream_s2mPipe_rData_twiceMode <= controlStream_s2mPipe_payload_twiceMode;
    end
    if(controlStream_s2mPipe_m2sPipe_ready) begin
      controlStream_s2mPipe_m2sPipe_rData_frameStart <= controlStream_s2mPipe_m2sPipe_payload_frameStart;
      controlStream_s2mPipe_m2sPipe_rData_rowEnd <= controlStream_s2mPipe_m2sPipe_payload_rowEnd;
      controlStream_s2mPipe_m2sPipe_rData_passMode <= controlStream_s2mPipe_m2sPipe_payload_passMode;
      controlStream_s2mPipe_m2sPipe_rData_passValid <= controlStream_s2mPipe_m2sPipe_payload_passValid;
      controlStream_s2mPipe_m2sPipe_rData_onceMode <= controlStream_s2mPipe_m2sPipe_payload_onceMode;
      controlStream_s2mPipe_m2sPipe_rData_onceValid <= controlStream_s2mPipe_m2sPipe_payload_onceValid;
      controlStream_s2mPipe_m2sPipe_rData_mainCompare <= controlStream_s2mPipe_m2sPipe_payload_mainCompare;
      controlStream_s2mPipe_m2sPipe_rData_counterCompare <= controlStream_s2mPipe_m2sPipe_payload_counterCompare;
      controlStream_s2mPipe_m2sPipe_rData_mainDiff <= controlStream_s2mPipe_m2sPipe_payload_mainDiff;
      controlStream_s2mPipe_m2sPipe_rData_counterDiff <= controlStream_s2mPipe_m2sPipe_payload_counterDiff;
      controlStream_s2mPipe_m2sPipe_rData_twiceCompValid <= controlStream_s2mPipe_m2sPipe_payload_twiceCompValid;
      controlStream_s2mPipe_m2sPipe_rData_twiceMode <= controlStream_s2mPipe_m2sPipe_payload_twiceMode;
    end
    if(controlStream_s2mPipe_m2sPipe_m2sPipe_ready) begin
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_frameStart <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_frameStart;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_rowEnd <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_rowEnd;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_passMode <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passMode;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_passValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_onceMode <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceMode;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_onceValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_twiceCompValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceCompValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_twiceMode <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceMode;
    end
    if(controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready) begin
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_frameStart <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_frameStart;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_rowEnd <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_rowEnd;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_passMode <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_passMode;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_passValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_passValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_onceMode <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_onceMode;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_onceValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_onceValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_twiceCompValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_twiceCompValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_twiceMode <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_twiceMode;
    end
    if(readStage_mainOnePixelStream_ready) begin
      readStage_mainOnePixelStream_rData <= readStage_mainOnePixelStream_payload;
    end
    if(readStage_mainOnePixelStream_s2mPipe_ready) begin
      readStage_mainOnePixelStream_s2mPipe_rData <= readStage_mainOnePixelStream_s2mPipe_payload;
    end
    if(readStage_counterOnePixelStream_ready) begin
      readStage_counterOnePixelStream_rData <= readStage_counterOnePixelStream_payload;
    end
    if(readStage_counterOnePixelStream_s2mPipe_ready) begin
      readStage_counterOnePixelStream_s2mPipe_rData <= readStage_counterOnePixelStream_s2mPipe_payload;
    end
    if(readStage_mainTwoPixelStream_ready) begin
      readStage_mainTwoPixelStream_rData <= readStage_mainTwoPixelStream_payload;
    end
    if(readStage_mainTwoPixelStream_s2mPipe_ready) begin
      readStage_mainTwoPixelStream_s2mPipe_rData <= readStage_mainTwoPixelStream_s2mPipe_payload;
    end
    if(readStage_counterTwoPixelStream_ready) begin
      readStage_counterTwoPixelStream_rData <= readStage_counterTwoPixelStream_payload;
    end
    if(readStage_counterTwoPixelStream_s2mPipe_ready) begin
      readStage_counterTwoPixelStream_s2mPipe_rData <= readStage_counterTwoPixelStream_s2mPipe_payload;
    end
    if(readStage_controlPipe_translated_ready) begin
      readStage_controlPipe_translated_rData_frameStart <= readStage_controlPipe_translated_payload_frameStart;
      readStage_controlPipe_translated_rData_rowEnd <= readStage_controlPipe_translated_payload_rowEnd;
      readStage_controlPipe_translated_rData_passMode <= readStage_controlPipe_translated_payload_passMode;
      readStage_controlPipe_translated_rData_passValid <= readStage_controlPipe_translated_payload_passValid;
      readStage_controlPipe_translated_rData_onceMode <= readStage_controlPipe_translated_payload_onceMode;
      readStage_controlPipe_translated_rData_onceValid <= readStage_controlPipe_translated_payload_onceValid;
      readStage_controlPipe_translated_rData_mainCompare <= readStage_controlPipe_translated_payload_mainCompare;
      readStage_controlPipe_translated_rData_counterCompare <= readStage_controlPipe_translated_payload_counterCompare;
      readStage_controlPipe_translated_rData_mainDiff <= readStage_controlPipe_translated_payload_mainDiff;
      readStage_controlPipe_translated_rData_counterDiff <= readStage_controlPipe_translated_payload_counterDiff;
      readStage_controlPipe_translated_rData_twiceCompValid <= readStage_controlPipe_translated_payload_twiceCompValid;
      readStage_controlPipe_translated_rData_twiceMode <= readStage_controlPipe_translated_payload_twiceMode;
    end
    if(readStage_controlPipe_translated_s2mPipe_ready) begin
      readStage_controlPipe_translated_s2mPipe_rData_frameStart <= readStage_controlPipe_translated_s2mPipe_payload_frameStart;
      readStage_controlPipe_translated_s2mPipe_rData_rowEnd <= readStage_controlPipe_translated_s2mPipe_payload_rowEnd;
      readStage_controlPipe_translated_s2mPipe_rData_passMode <= readStage_controlPipe_translated_s2mPipe_payload_passMode;
      readStage_controlPipe_translated_s2mPipe_rData_passValid <= readStage_controlPipe_translated_s2mPipe_payload_passValid;
      readStage_controlPipe_translated_s2mPipe_rData_onceMode <= readStage_controlPipe_translated_s2mPipe_payload_onceMode;
      readStage_controlPipe_translated_s2mPipe_rData_onceValid <= readStage_controlPipe_translated_s2mPipe_payload_onceValid;
      readStage_controlPipe_translated_s2mPipe_rData_mainCompare <= readStage_controlPipe_translated_s2mPipe_payload_mainCompare;
      readStage_controlPipe_translated_s2mPipe_rData_counterCompare <= readStage_controlPipe_translated_s2mPipe_payload_counterCompare;
      readStage_controlPipe_translated_s2mPipe_rData_mainDiff <= readStage_controlPipe_translated_s2mPipe_payload_mainDiff;
      readStage_controlPipe_translated_s2mPipe_rData_counterDiff <= readStage_controlPipe_translated_s2mPipe_payload_counterDiff;
      readStage_controlPipe_translated_s2mPipe_rData_twiceCompValid <= readStage_controlPipe_translated_s2mPipe_payload_twiceCompValid;
      readStage_controlPipe_translated_s2mPipe_rData_twiceMode <= readStage_controlPipe_translated_s2mPipe_payload_twiceMode;
    end
    if(compareStage_mainOnePixelStream_ready) begin
      compareStage_mainOnePixelStream_rData <= compareStage_mainOnePixelStream_payload;
    end
    if(compareStage_mainOnePixelStream_s2mPipe_ready) begin
      compareStage_mainOnePixelStream_s2mPipe_rData <= compareStage_mainOnePixelStream_s2mPipe_payload;
    end
    if(compareStage_counterOnePixelStream_ready) begin
      compareStage_counterOnePixelStream_rData <= compareStage_counterOnePixelStream_payload;
    end
    if(compareStage_counterOnePixelStream_s2mPipe_ready) begin
      compareStage_counterOnePixelStream_s2mPipe_rData <= compareStage_counterOnePixelStream_s2mPipe_payload;
    end
    if(compareStage_mainTwoPixelStream_ready) begin
      compareStage_mainTwoPixelStream_rData <= compareStage_mainTwoPixelStream_payload;
    end
    if(compareStage_mainTwoPixelStream_s2mPipe_ready) begin
      compareStage_mainTwoPixelStream_s2mPipe_rData <= compareStage_mainTwoPixelStream_s2mPipe_payload;
    end
    if(compareStage_counterTwoPixelStream_ready) begin
      compareStage_counterTwoPixelStream_rData <= compareStage_counterTwoPixelStream_payload;
    end
    if(compareStage_counterTwoPixelStream_s2mPipe_ready) begin
      compareStage_counterTwoPixelStream_s2mPipe_rData <= compareStage_counterTwoPixelStream_s2mPipe_payload;
    end
    if(compareStage_controlPipe_translated_ready) begin
      compareStage_controlPipe_translated_rData_frameStart <= compareStage_controlPipe_translated_payload_frameStart;
      compareStage_controlPipe_translated_rData_rowEnd <= compareStage_controlPipe_translated_payload_rowEnd;
      compareStage_controlPipe_translated_rData_passMode <= compareStage_controlPipe_translated_payload_passMode;
      compareStage_controlPipe_translated_rData_passValid <= compareStage_controlPipe_translated_payload_passValid;
      compareStage_controlPipe_translated_rData_onceMode <= compareStage_controlPipe_translated_payload_onceMode;
      compareStage_controlPipe_translated_rData_onceValid <= compareStage_controlPipe_translated_payload_onceValid;
      compareStage_controlPipe_translated_rData_mainCompare <= compareStage_controlPipe_translated_payload_mainCompare;
      compareStage_controlPipe_translated_rData_counterCompare <= compareStage_controlPipe_translated_payload_counterCompare;
      compareStage_controlPipe_translated_rData_mainDiff <= compareStage_controlPipe_translated_payload_mainDiff;
      compareStage_controlPipe_translated_rData_counterDiff <= compareStage_controlPipe_translated_payload_counterDiff;
      compareStage_controlPipe_translated_rData_twiceCompValid <= compareStage_controlPipe_translated_payload_twiceCompValid;
      compareStage_controlPipe_translated_rData_twiceMode <= compareStage_controlPipe_translated_payload_twiceMode;
    end
    if(compareStage_controlPipe_translated_s2mPipe_ready) begin
      compareStage_controlPipe_translated_s2mPipe_rData_frameStart <= compareStage_controlPipe_translated_s2mPipe_payload_frameStart;
      compareStage_controlPipe_translated_s2mPipe_rData_rowEnd <= compareStage_controlPipe_translated_s2mPipe_payload_rowEnd;
      compareStage_controlPipe_translated_s2mPipe_rData_passMode <= compareStage_controlPipe_translated_s2mPipe_payload_passMode;
      compareStage_controlPipe_translated_s2mPipe_rData_passValid <= compareStage_controlPipe_translated_s2mPipe_payload_passValid;
      compareStage_controlPipe_translated_s2mPipe_rData_onceMode <= compareStage_controlPipe_translated_s2mPipe_payload_onceMode;
      compareStage_controlPipe_translated_s2mPipe_rData_onceValid <= compareStage_controlPipe_translated_s2mPipe_payload_onceValid;
      compareStage_controlPipe_translated_s2mPipe_rData_mainCompare <= compareStage_controlPipe_translated_s2mPipe_payload_mainCompare;
      compareStage_controlPipe_translated_s2mPipe_rData_counterCompare <= compareStage_controlPipe_translated_s2mPipe_payload_counterCompare;
      compareStage_controlPipe_translated_s2mPipe_rData_mainDiff <= compareStage_controlPipe_translated_s2mPipe_payload_mainDiff;
      compareStage_controlPipe_translated_s2mPipe_rData_counterDiff <= compareStage_controlPipe_translated_s2mPipe_payload_counterDiff;
      compareStage_controlPipe_translated_s2mPipe_rData_twiceCompValid <= compareStage_controlPipe_translated_s2mPipe_payload_twiceCompValid;
      compareStage_controlPipe_translated_s2mPipe_rData_twiceMode <= compareStage_controlPipe_translated_s2mPipe_payload_twiceMode;
    end
    if(diffStage_mainOnePixelStream_ready) begin
      diffStage_mainOnePixelStream_rData <= diffStage_mainOnePixelStream_payload;
    end
    if(diffStage_mainOnePixelStream_s2mPipe_ready) begin
      diffStage_mainOnePixelStream_s2mPipe_rData <= diffStage_mainOnePixelStream_s2mPipe_payload;
    end
    if(diffStage_counterOnePixelStream_ready) begin
      diffStage_counterOnePixelStream_rData <= diffStage_counterOnePixelStream_payload;
    end
    if(diffStage_counterOnePixelStream_s2mPipe_ready) begin
      diffStage_counterOnePixelStream_s2mPipe_rData <= diffStage_counterOnePixelStream_s2mPipe_payload;
    end
    if(diffStage_mainTwoPixelStream_ready) begin
      diffStage_mainTwoPixelStream_rData <= diffStage_mainTwoPixelStream_payload;
    end
    if(diffStage_mainTwoPixelStream_s2mPipe_ready) begin
      diffStage_mainTwoPixelStream_s2mPipe_rData <= diffStage_mainTwoPixelStream_s2mPipe_payload;
    end
    if(diffStage_counterTwoPixelStream_ready) begin
      diffStage_counterTwoPixelStream_rData <= diffStage_counterTwoPixelStream_payload;
    end
    if(diffStage_counterTwoPixelStream_s2mPipe_ready) begin
      diffStage_counterTwoPixelStream_s2mPipe_rData <= diffStage_counterTwoPixelStream_s2mPipe_payload;
    end
    if(diffStage_controlPipe_fork_io_outputs_0_ready) begin
      diffStage_controlPipe_fork_io_outputs_0_rData_frameStart <= diffStage_controlPipe_fork_io_outputs_0_payload_frameStart;
      diffStage_controlPipe_fork_io_outputs_0_rData_rowEnd <= diffStage_controlPipe_fork_io_outputs_0_payload_rowEnd;
      diffStage_controlPipe_fork_io_outputs_0_rData_passMode <= diffStage_controlPipe_fork_io_outputs_0_payload_passMode;
      diffStage_controlPipe_fork_io_outputs_0_rData_passValid <= diffStage_controlPipe_fork_io_outputs_0_payload_passValid;
      diffStage_controlPipe_fork_io_outputs_0_rData_onceMode <= diffStage_controlPipe_fork_io_outputs_0_payload_onceMode;
      diffStage_controlPipe_fork_io_outputs_0_rData_onceValid <= diffStage_controlPipe_fork_io_outputs_0_payload_onceValid;
      diffStage_controlPipe_fork_io_outputs_0_rData_mainCompare <= diffStage_controlPipe_fork_io_outputs_0_payload_mainCompare;
      diffStage_controlPipe_fork_io_outputs_0_rData_counterCompare <= diffStage_controlPipe_fork_io_outputs_0_payload_counterCompare;
      diffStage_controlPipe_fork_io_outputs_0_rData_mainDiff <= diffStage_controlPipe_fork_io_outputs_0_payload_mainDiff;
      diffStage_controlPipe_fork_io_outputs_0_rData_counterDiff <= diffStage_controlPipe_fork_io_outputs_0_payload_counterDiff;
      diffStage_controlPipe_fork_io_outputs_0_rData_twiceCompValid <= diffStage_controlPipe_fork_io_outputs_0_payload_twiceCompValid;
      diffStage_controlPipe_fork_io_outputs_0_rData_twiceMode <= diffStage_controlPipe_fork_io_outputs_0_payload_twiceMode;
    end
    if(diffStage_controlPipe_fork_io_outputs_0_s2mPipe_ready) begin
      diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_frameStart <= diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_frameStart;
      diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_rowEnd <= diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_rowEnd;
      diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_passMode <= diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_passMode;
      diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_passValid <= diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_passValid;
      diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_onceMode <= diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_onceMode;
      diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_onceValid <= diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_onceValid;
      diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_mainCompare <= diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_mainCompare;
      diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_counterCompare <= diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_counterCompare;
      diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_mainDiff <= diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_mainDiff;
      diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_counterDiff <= diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_counterDiff;
      diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_twiceCompValid <= diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_twiceCompValid;
      diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_twiceMode <= diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_twiceMode;
    end
    if(resultStage_pixelStream_ready) begin
      resultStage_pixelStream_rData <= resultStage_pixelStream_payload;
    end
    if(resultStage_pixelStream_s2mPipe_ready) begin
      resultStage_pixelStream_s2mPipe_rData <= resultStage_pixelStream_s2mPipe_payload;
    end
    if(pixelsStream_ready) begin
      pixelsStream_rData_pixel <= pixelsStream_payload_pixel;
      pixelsStream_rData_frameStart <= pixelsStream_payload_frameStart;
      pixelsStream_rData_rowEnd <= pixelsStream_payload_rowEnd;
    end
    if(pixelsStream_s2mPipe_ready) begin
      pixelsStream_s2mPipe_rData_pixel <= pixelsStream_s2mPipe_payload_pixel;
      pixelsStream_s2mPipe_rData_frameStart <= pixelsStream_s2mPipe_payload_frameStart;
      pixelsStream_s2mPipe_rData_rowEnd <= pixelsStream_s2mPipe_payload_rowEnd;
    end
    if(pixelsIn_ready) begin
      pixelsIn_rData_pixel <= pixelsIn_payload_pixel;
      pixelsIn_rData_frameStart <= pixelsIn_payload_frameStart;
      pixelsIn_rData_rowEnd <= pixelsIn_payload_rowEnd;
    end
    if(pixelsIn_s2mPipe_ready) begin
      pixelsIn_s2mPipe_rData_pixel <= pixelsIn_s2mPipe_payload_pixel;
      pixelsIn_s2mPipe_rData_frameStart <= pixelsIn_s2mPipe_payload_frameStart;
      pixelsIn_s2mPipe_rData_rowEnd <= pixelsIn_s2mPipe_payload_rowEnd;
    end
  end


endmodule

module SuperResolutionPart3 (
  input               pixelsIn_valid,
  output reg          pixelsIn_ready,
  input      [7:0]    pixelsIn_payload_pixel,
  input               pixelsIn_payload_frameStart,
  input               pixelsIn_payload_rowEnd,
  input               pixelsIn_payload_inpValid,
  input               startIn,
  output reg          pixelsOut_valid,
  input               pixelsOut_ready,
  output reg [7:0]    pixelsOut_payload_pixel,
  output reg          pixelsOut_payload_frameStart,
  output reg          pixelsOut_payload_rowEnd,
  output reg          inpThreeDoneOut,
  input      [7:0]    thresholdIn,
  input      [9:0]    widthIn,
  input      [9:0]    heightIn,
  input               clk,
  input               resetn
);
  localparam controlStateMachine_enumDef_2_BOOT = 2'd0;
  localparam controlStateMachine_enumDef_2_HOLD = 2'd1;
  localparam controlStateMachine_enumDef_2_PASS = 2'd2;
  localparam controlStateMachine_enumDef_2_EXTRA = 2'd3;

  reg        [7:0]    CICC1851_lineBufferOne_port1;
  reg        [7:0]    CICC1851_lineBufferOne_port2;
  reg        [7:0]    CICC1851_lineBufferTwo_port1;
  reg        [7:0]    CICC1851_lineBufferTwo_port2;
  reg        [7:0]    CICC1851_lineBufferThree_port1;
  reg        [7:0]    CICC1851_lineBufferThree_port2;
  reg        [0:0]    CICC1851_validBufferOne_port1;
  reg        [0:0]    CICC1851_validBufferOne_port2;
  reg        [0:0]    CICC1851_validBufferTwo_port1;
  reg        [0:0]    CICC1851_validBufferTwo_port2;
  reg        [0:0]    CICC1851_validBufferThree_port1;
  reg        [0:0]    CICC1851_validBufferThree_port2;
  wire                diffStage_controlPipe_fork_io_input_ready;
  wire                diffStage_controlPipe_fork_io_outputs_0_valid;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_frameStart;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_rowEnd;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_pipeValid;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_firstRow;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_lastRow;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_finalResult;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_mainCompare;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_counterCompare;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_horizontalCompare;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_verticalCompare;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_payload_mainDiff;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_payload_counterDiff;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_payload_horizontalDiff;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_payload_verticalDiff;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_isHorizontalMin;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_payload_minDiff;
  wire       [1:0]    diffStage_controlPipe_fork_io_outputs_0_payload_currentPosition;
  wire       [1:0]    diffStage_controlPipe_fork_io_outputs_0_payload_nextPosition;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_horizontalDirectionValid;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_verticalDirectionValid;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_mainDirectionValid;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_counterDirectionValid;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_inValidMinDiff;
  wire                diffStage_controlPipe_fork_io_outputs_1_valid;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_frameStart;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_rowEnd;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_pipeValid;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_firstRow;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_lastRow;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_finalResult;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_mainCompare;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_counterCompare;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_horizontalCompare;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_verticalCompare;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_1_payload_horizontalDiff;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_1_payload_verticalDiff;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_isHorizontalMin;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_1_payload_minDiff;
  wire       [1:0]    diffStage_controlPipe_fork_io_outputs_1_payload_currentPosition;
  wire       [1:0]    diffStage_controlPipe_fork_io_outputs_1_payload_nextPosition;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_horizontalDirectionValid;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_verticalDirectionValid;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_mainDirectionValid;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_counterDirectionValid;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_inValidMinDiff;
  wire       [11:0]   CICC1851_bufferRowCount_valueNext;
  wire       [0:0]    CICC1851_bufferRowCount_valueNext_1;
  wire       [11:0]   CICC1851_bufferWAddr_valueNext;
  wire       [0:0]    CICC1851_bufferWAddr_valueNext_1;
  wire       [11:0]   CICC1851_outPixelAddr_valueNext;
  wire       [0:0]    CICC1851_outPixelAddr_valueNext_1;
  wire       [11:0]   CICC1851_outRowCount_valueNext;
  wire       [0:0]    CICC1851_outRowCount_valueNext_1;
  wire       [11:0]   CICC1851_alreadySendRow_valueNext;
  wire       [0:0]    CICC1851_alreadySendRow_valueNext_1;
  wire       [11:0]   CICC1851_alreadySendCountInRow_valueNext;
  wire       [0:0]    CICC1851_alreadySendCountInRow_valueNext_1;
  wire       [0:0]    CICC1851_nextRowBuffer;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l226;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l226_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l226_2;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l227;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l227_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l227_2;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l270;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l270_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l270_2;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l271;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l271_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l271_2;
  wire       [7:0]    CICC1851_lineBufferOne_port;
  wire                CICC1851_lineBufferOne_port_1;
  wire       [7:0]    CICC1851_lineBufferTwo_port;
  wire                CICC1851_lineBufferTwo_port_1;
  wire       [7:0]    CICC1851_lineBufferThree_port;
  wire                CICC1851_lineBufferThree_port_1;
  wire       [0:0]    CICC1851_validBufferOne_port;
  wire                CICC1851_validBufferOne_port_1;
  wire       [0:0]    CICC1851_validBufferTwo_port;
  wire                CICC1851_validBufferTwo_port_1;
  wire       [0:0]    CICC1851_validBufferThree_port;
  wire                CICC1851_validBufferThree_port_1;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_1;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_2;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_3;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_4;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_5;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_6;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_7;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_8;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_9;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_10;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_11;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_12;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_13;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_14;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_15;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_16;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_17;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_18;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_19;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_20;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_21;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_22;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_23;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_24;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_25;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_26;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_27;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_28;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_29;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_30;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_31;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_32;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_33;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_34;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_35;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_36;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_37;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_38;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_39;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_40;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_41;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_42;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_43;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_44;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_45;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_46;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_47;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_48;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_49;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_50;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_51;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_52;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_53;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_54;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_55;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_56;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_57;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_58;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_59;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_60;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_61;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_62;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_63;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_64;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_65;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_66;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_67;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_68;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_69;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_70;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_71;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_72;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_73;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_74;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_75;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_76;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_77;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_78;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_79;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_80;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_81;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_82;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_83;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_84;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_85;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_86;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_87;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_88;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_89;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_90;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_91;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_92;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_93;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_94;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_95;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_96;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_97;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_98;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_99;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_100;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_101;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_102;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_103;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_104;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_105;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_106;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_107;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_108;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_109;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_110;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_111;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_112;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_113;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_114;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_115;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_116;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_117;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_118;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_119;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_120;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_121;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_122;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_123;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_124;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_125;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_126;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_127;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_128;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_129;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_130;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_131;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_132;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_133;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_134;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_135;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_136;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_137;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_138;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_139;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_140;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_141;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_142;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_143;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_144;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_145;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_146;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_147;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_148;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_149;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_150;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_151;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_152;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_153;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_154;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_155;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_156;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_157;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_158;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_159;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_160;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_161;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_162;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_163;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_164;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_165;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_166;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_167;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_168;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_169;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_170;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_171;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_172;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_173;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_174;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_175;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_176;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_177;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_178;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_179;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_180;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_181;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_182;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_183;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_184;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_185;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_186;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_187;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_188;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_189;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_190;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_191;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_192;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_193;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_194;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_195;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_196;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_197;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_198;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_199;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_200;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_201;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_202;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_203;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_204;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_205;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_206;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_207;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_208;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_209;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_210;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_211;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_212;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_213;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_214;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_215;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_216;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_217;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_218;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_219;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_220;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_221;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_222;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_223;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_224;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_225;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_226;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_227;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_228;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_229;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_230;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_231;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_232;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_233;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_234;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_235;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_236;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_237;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_238;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_239;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_240;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_241;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_242;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_243;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_244;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_245;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_246;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_247;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_248;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_249;
  wire       [11:0]   CICC1851_when_SuperResolutionPart3_l1202;
  wire       [11:0]   CICC1851_when_SuperResolutionPart3_l1205;
  wire       [11:0]   CICC1851_when_SuperResolutionPart3_l1205_1;
  wire       [11:0]   CICC1851_when_SuperResolutionPart3_l1205_2;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l1223;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l1223_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l1223_2;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l1224;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l1224_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart3_l1224_2;
  reg                 inpThreeDone;
  reg                 startIn_regNext;
  wire                when_SuperResolutionPart3_l72;
  reg                 readDone;
  wire                when_SuperResolutionPart3_l75;
  reg                 startRead;
  wire                when_SuperResolutionPart3_l78;
  wire                when_SuperResolutionPart3_l78_1;
  reg                 frameStart;
  reg        [7:0]    inpThreshold;
  reg        [9:0]    bmpWidth;
  reg        [9:0]    bmpHeight;
  reg                 holdBuffer;
  wire                when_SuperResolutionPart3_l93;
  reg                 writeDone;
  wire                when_SuperResolutionPart3_l96;
  reg                 bufferRowCount_willIncrement;
  reg                 bufferRowCount_willClear;
  reg        [11:0]   bufferRowCount_valueNext;
  reg        [11:0]   bufferRowCount_value;
  wire                bufferRowCount_willOverflowIfInc;
  wire                bufferRowCount_willOverflow;
  reg                 bufferEnable;
  wire                when_SuperResolutionPart3_l102;
  wire                when_SuperResolutionPart3_l102_1;
  reg        [1:0]    bufferSwitch;
  reg        [1:0]    nextRowBuffer;
  reg        [1:0]    currentRowBuffer;
  reg                 bufferReuse;
  reg                 bufferWAddr_willIncrement;
  reg                 bufferWAddr_willClear;
  reg        [11:0]   bufferWAddr_valueNext;
  reg        [11:0]   bufferWAddr_value;
  wire                bufferWAddr_willOverflowIfInc;
  wire                bufferWAddr_willOverflow;
  reg                 outPixelAddr_willIncrement;
  reg                 outPixelAddr_willClear;
  reg        [11:0]   outPixelAddr_valueNext;
  reg        [11:0]   outPixelAddr_value;
  wire                outPixelAddr_willOverflowIfInc;
  wire                outPixelAddr_willOverflow;
  reg                 outRowCount_willIncrement;
  reg                 outRowCount_willClear;
  reg        [11:0]   outRowCount_valueNext;
  reg        [11:0]   outRowCount_value;
  wire                outRowCount_willOverflowIfInc;
  wire                outRowCount_willOverflow;
  reg                 alreadySendRow_willIncrement;
  reg                 alreadySendRow_willClear;
  reg        [11:0]   alreadySendRow_valueNext;
  reg        [11:0]   alreadySendRow_value;
  wire                alreadySendRow_willOverflowIfInc;
  wire                alreadySendRow_willOverflow;
  reg                 alreadySendCountInRow_willIncrement;
  reg                 alreadySendCountInRow_willClear;
  reg        [11:0]   alreadySendCountInRow_valueNext;
  reg        [11:0]   alreadySendCountInRow_value;
  wire                alreadySendCountInRow_willOverflowIfInc;
  wire                alreadySendCountInRow_willOverflow;
  reg                 alreadyReachRowEnd;
  reg                 alreadyReachFinalRow;
  reg                 outReachRowEnd;
  reg                 outReachFinalRow;
  reg                 bufferReachRowEnd;
  reg                 bufferReachFinalRow;
  reg        [7:0]    minDiff;
  reg        [7:0]    candidatePixel;
  reg                 isHorizontalDirection;
  reg                 inValidMinDiff;
  reg                 startIn_regNext_1;
  wire                when_SuperResolutionPart3_l154;
  reg        [11:0]   mainAddrOne;
  reg        [11:0]   counterAddrOne;
  reg        [11:0]   mainAddrTwo;
  reg        [11:0]   counterAddrTwo;
  reg        [11:0]   mainAddrThree;
  reg        [11:0]   counterAddrThree;
  wire                validStream_valid;
  reg                 validStream_ready;
  wire                controlStream_valid;
  wire                controlStream_ready;
  wire                controlStream_payload_frameStart;
  wire                controlStream_payload_rowEnd;
  wire                controlStream_payload_pipeValid;
  wire                controlStream_payload_firstRow;
  wire                controlStream_payload_lastRow;
  wire                controlStream_payload_finalResult;
  wire                controlStream_payload_mainCompare;
  wire                controlStream_payload_counterCompare;
  wire                controlStream_payload_horizontalCompare;
  wire                controlStream_payload_verticalCompare;
  wire       [7:0]    controlStream_payload_mainDiff;
  wire       [7:0]    controlStream_payload_counterDiff;
  wire       [7:0]    controlStream_payload_horizontalDiff;
  wire       [7:0]    controlStream_payload_verticalDiff;
  wire                controlStream_payload_isHorizontalMin;
  wire       [7:0]    controlStream_payload_minDiff;
  wire       [1:0]    controlStream_payload_currentPosition;
  wire       [1:0]    controlStream_payload_nextPosition;
  wire                controlStream_payload_horizontalDirectionValid;
  wire                controlStream_payload_verticalDirectionValid;
  wire                controlStream_payload_mainDirectionValid;
  wire                controlStream_payload_counterDirectionValid;
  wire                controlStream_payload_inValidMinDiff;
  reg                 controls_frameStart;
  reg                 controls_rowEnd;
  reg                 controls_pipeValid;
  reg                 controls_firstRow;
  reg                 controls_lastRow;
  reg                 controls_finalResult;
  wire                controls_mainCompare;
  wire                controls_counterCompare;
  wire                controls_horizontalCompare;
  wire                controls_verticalCompare;
  wire       [7:0]    controls_mainDiff;
  wire       [7:0]    controls_counterDiff;
  wire       [7:0]    controls_horizontalDiff;
  wire       [7:0]    controls_verticalDiff;
  wire                controls_isHorizontalMin;
  wire       [7:0]    controls_minDiff;
  reg        [1:0]    controls_currentPosition;
  reg        [1:0]    controls_nextPosition;
  wire                controls_horizontalDirectionValid;
  wire                controls_verticalDirectionValid;
  wire                controls_mainDirectionValid;
  wire                controls_counterDirectionValid;
  wire                controls_inValidMinDiff;
  wire       [59:0]   CICC1851_controls_frameStart;
  wire                mainPixelAddrOneStream_valid;
  wire                mainPixelAddrOneStream_ready;
  wire       [11:0]   mainPixelAddrOneStream_payload;
  wire                counterPixelAddrOneStream_valid;
  wire                counterPixelAddrOneStream_ready;
  wire       [11:0]   counterPixelAddrOneStream_payload;
  wire                mainPixelAddrTwoStream_valid;
  wire                mainPixelAddrTwoStream_ready;
  wire       [11:0]   mainPixelAddrTwoStream_payload;
  wire                counterPixelAddrTwoStream_valid;
  wire                counterPixelAddrTwoStream_ready;
  wire       [11:0]   counterPixelAddrTwoStream_payload;
  wire                mainPixelAddrThreeStream_valid;
  wire                mainPixelAddrThreeStream_ready;
  wire       [11:0]   mainPixelAddrThreeStream_payload;
  wire                counterPixelAddrThreeStream_valid;
  wire                counterPixelAddrThreeStream_ready;
  wire       [11:0]   counterPixelAddrThreeStream_payload;
  wire                mainValidAddrOneStream_valid;
  wire                mainValidAddrOneStream_ready;
  wire       [11:0]   mainValidAddrOneStream_payload;
  wire                counterValidAddrOneStream_valid;
  wire                counterValidAddrOneStream_ready;
  wire       [11:0]   counterValidAddrOneStream_payload;
  wire                mainValidAddrTwoStream_valid;
  wire                mainValidAddrTwoStream_ready;
  wire       [11:0]   mainValidAddrTwoStream_payload;
  wire                counterValidAddrTwoStream_valid;
  wire                counterValidAddrTwoStream_ready;
  wire       [11:0]   counterValidAddrTwoStream_payload;
  wire                mainValidAddrThreeStream_valid;
  wire                mainValidAddrThreeStream_ready;
  wire       [11:0]   mainValidAddrThreeStream_payload;
  wire                counterValidAddrThreeStream_valid;
  wire                counterValidAddrThreeStream_ready;
  wire       [11:0]   counterValidAddrThreeStream_payload;
  wire                pixelsIn_s2mPipe_valid;
  reg                 pixelsIn_s2mPipe_ready;
  wire       [7:0]    pixelsIn_s2mPipe_payload_pixel;
  wire                pixelsIn_s2mPipe_payload_frameStart;
  wire                pixelsIn_s2mPipe_payload_rowEnd;
  wire                pixelsIn_s2mPipe_payload_inpValid;
  reg                 pixelsIn_rValid;
  reg        [7:0]    pixelsIn_rData_pixel;
  reg                 pixelsIn_rData_frameStart;
  reg                 pixelsIn_rData_rowEnd;
  reg                 pixelsIn_rData_inpValid;
  wire                pixelsIn_s2mPipe_m2sPipe_valid;
  wire                pixelsIn_s2mPipe_m2sPipe_ready;
  wire       [7:0]    pixelsIn_s2mPipe_m2sPipe_payload_pixel;
  wire                pixelsIn_s2mPipe_m2sPipe_payload_frameStart;
  wire                pixelsIn_s2mPipe_m2sPipe_payload_rowEnd;
  wire                pixelsIn_s2mPipe_m2sPipe_payload_inpValid;
  reg                 pixelsIn_s2mPipe_rValid;
  reg        [7:0]    pixelsIn_s2mPipe_rData_pixel;
  reg                 pixelsIn_s2mPipe_rData_frameStart;
  reg                 pixelsIn_s2mPipe_rData_rowEnd;
  reg                 pixelsIn_s2mPipe_rData_inpValid;
  wire                when_Stream_l368;
  wire                passPixels_valid;
  wire                passPixels_ready;
  wire       [7:0]    passPixels_payload_pixel;
  wire                passPixels_payload_frameStart;
  wire                passPixels_payload_rowEnd;
  wire                passPixels_payload_inpValid;
  wire                passPixels_fire;
  wire                when_SuperResolutionPart3_l226;
  wire                passPixels_fire_1;
  wire                when_SuperResolutionPart3_l227;
  wire                passPixels_fire_2;
  wire                when_SuperResolutionPart3_l230;
  wire                passPixels_fire_3;
  wire                when_SuperResolutionPart3_l243;
  wire                when_SuperResolutionPart3_l244;
  wire                passPixels_fire_4;
  wire                when_SuperResolutionPart3_l251;
  wire                when_SuperResolutionPart3_l255;
  wire                passPixels_fire_5;
  wire                when_SuperResolutionPart3_l262;
  wire                pixelsOut_fire;
  wire                when_SuperResolutionPart3_l270;
  wire                pixelsOut_fire_1;
  wire                when_SuperResolutionPart3_l271;
  wire                pixelsOut_fire_2;
  wire                pixelsOut_fire_3;
  wire                when_SuperResolutionPart3_l282;
  wire                passPixels_fire_6;
  wire                passPixels_fire_7;
  wire                passPixels_fire_8;
  wire                passPixels_fire_9;
  wire                passPixels_fire_10;
  wire                passPixels_fire_11;
  wire                passPixels_fire_12;
  wire                mainPixelAddrOneStream_s2mPipe_valid;
  reg                 mainPixelAddrOneStream_s2mPipe_ready;
  wire       [11:0]   mainPixelAddrOneStream_s2mPipe_payload;
  reg                 mainPixelAddrOneStream_rValid;
  reg        [11:0]   mainPixelAddrOneStream_rData;
  wire                mainPixelAddrOneStream_s2mPipe_m2sPipe_valid;
  wire                mainPixelAddrOneStream_s2mPipe_m2sPipe_ready;
  wire       [11:0]   mainPixelAddrOneStream_s2mPipe_m2sPipe_payload;
  reg                 mainPixelAddrOneStream_s2mPipe_rValid;
  reg        [11:0]   mainPixelAddrOneStream_s2mPipe_rData;
  wire                when_Stream_l368_1;
  wire                CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_mainOnePixelStream_payload;
  reg                 CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_1;
  reg                 CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_mainOnePixelStream_payload_1;
  wire                readStage_mainOnePixelStream_valid;
  wire                readStage_mainOnePixelStream_ready;
  wire       [7:0]    readStage_mainOnePixelStream_payload;
  reg                 CICC1851_readStage_mainOnePixelStream_valid;
  reg        [7:0]    CICC1851_readStage_mainOnePixelStream_payload_2;
  wire                when_Stream_l368_2;
  wire                counterPixelAddrOneStream_s2mPipe_valid;
  reg                 counterPixelAddrOneStream_s2mPipe_ready;
  wire       [11:0]   counterPixelAddrOneStream_s2mPipe_payload;
  reg                 counterPixelAddrOneStream_rValid;
  reg        [11:0]   counterPixelAddrOneStream_rData;
  wire                counterPixelAddrOneStream_s2mPipe_m2sPipe_valid;
  wire                counterPixelAddrOneStream_s2mPipe_m2sPipe_ready;
  wire       [11:0]   counterPixelAddrOneStream_s2mPipe_m2sPipe_payload;
  reg                 counterPixelAddrOneStream_s2mPipe_rValid;
  reg        [11:0]   counterPixelAddrOneStream_s2mPipe_rData;
  wire                when_Stream_l368_3;
  wire                CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_counterOnePixelStream_payload;
  reg                 CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_2;
  reg                 CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_counterOnePixelStream_payload_1;
  wire                readStage_counterOnePixelStream_valid;
  wire                readStage_counterOnePixelStream_ready;
  wire       [7:0]    readStage_counterOnePixelStream_payload;
  reg                 CICC1851_readStage_counterOnePixelStream_valid;
  reg        [7:0]    CICC1851_readStage_counterOnePixelStream_payload_2;
  wire                when_Stream_l368_4;
  wire                mainPixelAddrTwoStream_s2mPipe_valid;
  reg                 mainPixelAddrTwoStream_s2mPipe_ready;
  wire       [11:0]   mainPixelAddrTwoStream_s2mPipe_payload;
  reg                 mainPixelAddrTwoStream_rValid;
  reg        [11:0]   mainPixelAddrTwoStream_rData;
  wire                mainPixelAddrTwoStream_s2mPipe_m2sPipe_valid;
  wire                mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire       [11:0]   mainPixelAddrTwoStream_s2mPipe_m2sPipe_payload;
  reg                 mainPixelAddrTwoStream_s2mPipe_rValid;
  reg        [11:0]   mainPixelAddrTwoStream_s2mPipe_rData;
  wire                when_Stream_l368_5;
  wire                CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_mainTwoPixelStream_payload;
  reg                 CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_3;
  reg                 CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_mainTwoPixelStream_payload_1;
  wire                readStage_mainTwoPixelStream_valid;
  wire                readStage_mainTwoPixelStream_ready;
  wire       [7:0]    readStage_mainTwoPixelStream_payload;
  reg                 CICC1851_readStage_mainTwoPixelStream_valid;
  reg        [7:0]    CICC1851_readStage_mainTwoPixelStream_payload_2;
  wire                when_Stream_l368_6;
  wire                counterPixelAddrTwoStream_s2mPipe_valid;
  reg                 counterPixelAddrTwoStream_s2mPipe_ready;
  wire       [11:0]   counterPixelAddrTwoStream_s2mPipe_payload;
  reg                 counterPixelAddrTwoStream_rValid;
  reg        [11:0]   counterPixelAddrTwoStream_rData;
  wire                counterPixelAddrTwoStream_s2mPipe_m2sPipe_valid;
  wire                counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire       [11:0]   counterPixelAddrTwoStream_s2mPipe_m2sPipe_payload;
  reg                 counterPixelAddrTwoStream_s2mPipe_rValid;
  reg        [11:0]   counterPixelAddrTwoStream_s2mPipe_rData;
  wire                when_Stream_l368_7;
  wire                CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_counterTwoPixelStream_payload;
  reg                 CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_4;
  reg                 CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_counterTwoPixelStream_payload_1;
  wire                readStage_counterTwoPixelStream_valid;
  wire                readStage_counterTwoPixelStream_ready;
  wire       [7:0]    readStage_counterTwoPixelStream_payload;
  reg                 CICC1851_readStage_counterTwoPixelStream_valid;
  reg        [7:0]    CICC1851_readStage_counterTwoPixelStream_payload_2;
  wire                when_Stream_l368_8;
  wire                mainPixelAddrThreeStream_s2mPipe_valid;
  reg                 mainPixelAddrThreeStream_s2mPipe_ready;
  wire       [11:0]   mainPixelAddrThreeStream_s2mPipe_payload;
  reg                 mainPixelAddrThreeStream_rValid;
  reg        [11:0]   mainPixelAddrThreeStream_rData;
  wire                mainPixelAddrThreeStream_s2mPipe_m2sPipe_valid;
  wire                mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready;
  wire       [11:0]   mainPixelAddrThreeStream_s2mPipe_m2sPipe_payload;
  reg                 mainPixelAddrThreeStream_s2mPipe_rValid;
  reg        [11:0]   mainPixelAddrThreeStream_s2mPipe_rData;
  wire                when_Stream_l368_9;
  wire                CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_mainThreePixelStream_payload;
  reg                 CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_5;
  reg                 CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_mainThreePixelStream_payload_1;
  wire                readStage_mainThreePixelStream_valid;
  wire                readStage_mainThreePixelStream_ready;
  wire       [7:0]    readStage_mainThreePixelStream_payload;
  reg                 CICC1851_readStage_mainThreePixelStream_valid;
  reg        [7:0]    CICC1851_readStage_mainThreePixelStream_payload_2;
  wire                when_Stream_l368_10;
  wire                counterPixelAddrThreeStream_s2mPipe_valid;
  reg                 counterPixelAddrThreeStream_s2mPipe_ready;
  wire       [11:0]   counterPixelAddrThreeStream_s2mPipe_payload;
  reg                 counterPixelAddrThreeStream_rValid;
  reg        [11:0]   counterPixelAddrThreeStream_rData;
  wire                counterPixelAddrThreeStream_s2mPipe_m2sPipe_valid;
  wire                counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready;
  wire       [11:0]   counterPixelAddrThreeStream_s2mPipe_m2sPipe_payload;
  reg                 counterPixelAddrThreeStream_s2mPipe_rValid;
  reg        [11:0]   counterPixelAddrThreeStream_s2mPipe_rData;
  wire                when_Stream_l368_11;
  wire                CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_counterThreePixelStream_payload;
  reg                 CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_6;
  reg                 CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_counterThreePixelStream_payload_1;
  wire                readStage_counterThreePixelStream_valid;
  wire                readStage_counterThreePixelStream_ready;
  wire       [7:0]    readStage_counterThreePixelStream_payload;
  reg                 CICC1851_readStage_counterThreePixelStream_valid;
  reg        [7:0]    CICC1851_readStage_counterThreePixelStream_payload_2;
  wire                when_Stream_l368_12;
  wire                mainValidAddrOneStream_s2mPipe_valid;
  reg                 mainValidAddrOneStream_s2mPipe_ready;
  wire       [11:0]   mainValidAddrOneStream_s2mPipe_payload;
  reg                 mainValidAddrOneStream_rValid;
  reg        [11:0]   mainValidAddrOneStream_rData;
  wire                mainValidAddrOneStream_s2mPipe_m2sPipe_valid;
  wire                mainValidAddrOneStream_s2mPipe_m2sPipe_ready;
  wire       [11:0]   mainValidAddrOneStream_s2mPipe_m2sPipe_payload;
  reg                 mainValidAddrOneStream_s2mPipe_rValid;
  reg        [11:0]   mainValidAddrOneStream_s2mPipe_rData;
  wire                when_Stream_l368_13;
  wire                CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_1;
  wire                CICC1851_readStage_mainOneValidStream_payload;
  reg                 CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_7;
  reg                 CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_3;
  reg                 CICC1851_readStage_mainOneValidStream_payload_1;
  wire                readStage_mainOneValidStream_valid;
  wire                readStage_mainOneValidStream_ready;
  wire                readStage_mainOneValidStream_payload;
  reg                 CICC1851_readStage_mainOneValidStream_valid;
  reg                 CICC1851_readStage_mainOneValidStream_payload_2;
  wire                when_Stream_l368_14;
  wire                counterValidAddrOneStream_s2mPipe_valid;
  reg                 counterValidAddrOneStream_s2mPipe_ready;
  wire       [11:0]   counterValidAddrOneStream_s2mPipe_payload;
  reg                 counterValidAddrOneStream_rValid;
  reg        [11:0]   counterValidAddrOneStream_rData;
  wire                counterValidAddrOneStream_s2mPipe_m2sPipe_valid;
  wire                counterValidAddrOneStream_s2mPipe_m2sPipe_ready;
  wire       [11:0]   counterValidAddrOneStream_s2mPipe_m2sPipe_payload;
  reg                 counterValidAddrOneStream_s2mPipe_rValid;
  reg        [11:0]   counterValidAddrOneStream_s2mPipe_rData;
  wire                when_Stream_l368_15;
  wire                CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_1;
  wire                CICC1851_readStage_counterOneValidStream_payload;
  reg                 CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_8;
  reg                 CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_3;
  reg                 CICC1851_readStage_counterOneValidStream_payload_1;
  wire                readStage_counterOneValidStream_valid;
  wire                readStage_counterOneValidStream_ready;
  wire                readStage_counterOneValidStream_payload;
  reg                 CICC1851_readStage_counterOneValidStream_valid;
  reg                 CICC1851_readStage_counterOneValidStream_payload_2;
  wire                when_Stream_l368_16;
  wire                mainValidAddrTwoStream_s2mPipe_valid;
  reg                 mainValidAddrTwoStream_s2mPipe_ready;
  wire       [11:0]   mainValidAddrTwoStream_s2mPipe_payload;
  reg                 mainValidAddrTwoStream_rValid;
  reg        [11:0]   mainValidAddrTwoStream_rData;
  wire                mainValidAddrTwoStream_s2mPipe_m2sPipe_valid;
  wire                mainValidAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire       [11:0]   mainValidAddrTwoStream_s2mPipe_m2sPipe_payload;
  reg                 mainValidAddrTwoStream_s2mPipe_rValid;
  reg        [11:0]   mainValidAddrTwoStream_s2mPipe_rData;
  wire                when_Stream_l368_17;
  wire                CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_1;
  wire                CICC1851_readStage_mainTwoValidStream_payload;
  reg                 CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_9;
  reg                 CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_3;
  reg                 CICC1851_readStage_mainTwoValidStream_payload_1;
  wire                readStage_mainTwoValidStream_valid;
  wire                readStage_mainTwoValidStream_ready;
  wire                readStage_mainTwoValidStream_payload;
  reg                 CICC1851_readStage_mainTwoValidStream_valid;
  reg                 CICC1851_readStage_mainTwoValidStream_payload_2;
  wire                when_Stream_l368_18;
  wire                counterValidAddrTwoStream_s2mPipe_valid;
  reg                 counterValidAddrTwoStream_s2mPipe_ready;
  wire       [11:0]   counterValidAddrTwoStream_s2mPipe_payload;
  reg                 counterValidAddrTwoStream_rValid;
  reg        [11:0]   counterValidAddrTwoStream_rData;
  wire                counterValidAddrTwoStream_s2mPipe_m2sPipe_valid;
  wire                counterValidAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire       [11:0]   counterValidAddrTwoStream_s2mPipe_m2sPipe_payload;
  reg                 counterValidAddrTwoStream_s2mPipe_rValid;
  reg        [11:0]   counterValidAddrTwoStream_s2mPipe_rData;
  wire                when_Stream_l368_19;
  wire                CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_1;
  wire                CICC1851_readStage_counterTwoValidStream_payload;
  reg                 CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_10;
  reg                 CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_3;
  reg                 CICC1851_readStage_counterTwoValidStream_payload_1;
  wire                readStage_counterTwoValidStream_valid;
  wire                readStage_counterTwoValidStream_ready;
  wire                readStage_counterTwoValidStream_payload;
  reg                 CICC1851_readStage_counterTwoValidStream_valid;
  reg                 CICC1851_readStage_counterTwoValidStream_payload_2;
  wire                when_Stream_l368_20;
  wire                mainValidAddrThreeStream_s2mPipe_valid;
  reg                 mainValidAddrThreeStream_s2mPipe_ready;
  wire       [11:0]   mainValidAddrThreeStream_s2mPipe_payload;
  reg                 mainValidAddrThreeStream_rValid;
  reg        [11:0]   mainValidAddrThreeStream_rData;
  wire                mainValidAddrThreeStream_s2mPipe_m2sPipe_valid;
  wire                mainValidAddrThreeStream_s2mPipe_m2sPipe_ready;
  wire       [11:0]   mainValidAddrThreeStream_s2mPipe_m2sPipe_payload;
  reg                 mainValidAddrThreeStream_s2mPipe_rValid;
  reg        [11:0]   mainValidAddrThreeStream_s2mPipe_rData;
  wire                when_Stream_l368_21;
  wire                CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_1;
  wire                CICC1851_readStage_mainThreeValidStream_payload;
  reg                 CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_11;
  reg                 CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_3;
  reg                 CICC1851_readStage_mainThreeValidStream_payload_1;
  wire                readStage_mainThreeValidStream_valid;
  wire                readStage_mainThreeValidStream_ready;
  wire                readStage_mainThreeValidStream_payload;
  reg                 CICC1851_readStage_mainThreeValidStream_valid;
  reg                 CICC1851_readStage_mainThreeValidStream_payload_2;
  wire                when_Stream_l368_22;
  wire                counterValidAddrThreeStream_s2mPipe_valid;
  reg                 counterValidAddrThreeStream_s2mPipe_ready;
  wire       [11:0]   counterValidAddrThreeStream_s2mPipe_payload;
  reg                 counterValidAddrThreeStream_rValid;
  reg        [11:0]   counterValidAddrThreeStream_rData;
  wire                counterValidAddrThreeStream_s2mPipe_m2sPipe_valid;
  wire                counterValidAddrThreeStream_s2mPipe_m2sPipe_ready;
  wire       [11:0]   counterValidAddrThreeStream_s2mPipe_m2sPipe_payload;
  reg                 counterValidAddrThreeStream_s2mPipe_rValid;
  reg        [11:0]   counterValidAddrThreeStream_s2mPipe_rData;
  wire                when_Stream_l368_23;
  wire                CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_1;
  wire                CICC1851_readStage_counterThreeValidStream_payload;
  reg                 CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_12;
  reg                 CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_3;
  reg                 CICC1851_readStage_counterThreeValidStream_payload_1;
  wire                readStage_counterThreeValidStream_valid;
  wire                readStage_counterThreeValidStream_ready;
  wire                readStage_counterThreeValidStream_payload;
  reg                 CICC1851_readStage_counterThreeValidStream_valid;
  reg                 CICC1851_readStage_counterThreeValidStream_payload_2;
  wire                when_Stream_l368_24;
  wire                controlStream_s2mPipe_valid;
  reg                 controlStream_s2mPipe_ready;
  wire                controlStream_s2mPipe_payload_frameStart;
  wire                controlStream_s2mPipe_payload_rowEnd;
  wire                controlStream_s2mPipe_payload_pipeValid;
  wire                controlStream_s2mPipe_payload_firstRow;
  wire                controlStream_s2mPipe_payload_lastRow;
  wire                controlStream_s2mPipe_payload_finalResult;
  wire                controlStream_s2mPipe_payload_mainCompare;
  wire                controlStream_s2mPipe_payload_counterCompare;
  wire                controlStream_s2mPipe_payload_horizontalCompare;
  wire                controlStream_s2mPipe_payload_verticalCompare;
  wire       [7:0]    controlStream_s2mPipe_payload_mainDiff;
  wire       [7:0]    controlStream_s2mPipe_payload_counterDiff;
  wire       [7:0]    controlStream_s2mPipe_payload_horizontalDiff;
  wire       [7:0]    controlStream_s2mPipe_payload_verticalDiff;
  wire                controlStream_s2mPipe_payload_isHorizontalMin;
  wire       [7:0]    controlStream_s2mPipe_payload_minDiff;
  wire       [1:0]    controlStream_s2mPipe_payload_currentPosition;
  wire       [1:0]    controlStream_s2mPipe_payload_nextPosition;
  wire                controlStream_s2mPipe_payload_horizontalDirectionValid;
  wire                controlStream_s2mPipe_payload_verticalDirectionValid;
  wire                controlStream_s2mPipe_payload_mainDirectionValid;
  wire                controlStream_s2mPipe_payload_counterDirectionValid;
  wire                controlStream_s2mPipe_payload_inValidMinDiff;
  reg                 controlStream_rValid;
  reg                 controlStream_rData_frameStart;
  reg                 controlStream_rData_rowEnd;
  reg                 controlStream_rData_pipeValid;
  reg                 controlStream_rData_firstRow;
  reg                 controlStream_rData_lastRow;
  reg                 controlStream_rData_finalResult;
  reg                 controlStream_rData_mainCompare;
  reg                 controlStream_rData_counterCompare;
  reg                 controlStream_rData_horizontalCompare;
  reg                 controlStream_rData_verticalCompare;
  reg        [7:0]    controlStream_rData_mainDiff;
  reg        [7:0]    controlStream_rData_counterDiff;
  reg        [7:0]    controlStream_rData_horizontalDiff;
  reg        [7:0]    controlStream_rData_verticalDiff;
  reg                 controlStream_rData_isHorizontalMin;
  reg        [7:0]    controlStream_rData_minDiff;
  reg        [1:0]    controlStream_rData_currentPosition;
  reg        [1:0]    controlStream_rData_nextPosition;
  reg                 controlStream_rData_horizontalDirectionValid;
  reg                 controlStream_rData_verticalDirectionValid;
  reg                 controlStream_rData_mainDirectionValid;
  reg                 controlStream_rData_counterDirectionValid;
  reg                 controlStream_rData_inValidMinDiff;
  wire                controlStream_s2mPipe_m2sPipe_valid;
  reg                 controlStream_s2mPipe_m2sPipe_ready;
  wire                controlStream_s2mPipe_m2sPipe_payload_frameStart;
  wire                controlStream_s2mPipe_m2sPipe_payload_rowEnd;
  wire                controlStream_s2mPipe_m2sPipe_payload_pipeValid;
  wire                controlStream_s2mPipe_m2sPipe_payload_firstRow;
  wire                controlStream_s2mPipe_m2sPipe_payload_lastRow;
  wire                controlStream_s2mPipe_m2sPipe_payload_finalResult;
  wire                controlStream_s2mPipe_m2sPipe_payload_mainCompare;
  wire                controlStream_s2mPipe_m2sPipe_payload_counterCompare;
  wire                controlStream_s2mPipe_m2sPipe_payload_horizontalCompare;
  wire                controlStream_s2mPipe_m2sPipe_payload_verticalCompare;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_payload_mainDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_payload_counterDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_payload_horizontalDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_payload_verticalDiff;
  wire                controlStream_s2mPipe_m2sPipe_payload_isHorizontalMin;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_payload_minDiff;
  wire       [1:0]    controlStream_s2mPipe_m2sPipe_payload_currentPosition;
  wire       [1:0]    controlStream_s2mPipe_m2sPipe_payload_nextPosition;
  wire                controlStream_s2mPipe_m2sPipe_payload_horizontalDirectionValid;
  wire                controlStream_s2mPipe_m2sPipe_payload_verticalDirectionValid;
  wire                controlStream_s2mPipe_m2sPipe_payload_mainDirectionValid;
  wire                controlStream_s2mPipe_m2sPipe_payload_counterDirectionValid;
  wire                controlStream_s2mPipe_m2sPipe_payload_inValidMinDiff;
  reg                 controlStream_s2mPipe_rValid;
  reg                 controlStream_s2mPipe_rData_frameStart;
  reg                 controlStream_s2mPipe_rData_rowEnd;
  reg                 controlStream_s2mPipe_rData_pipeValid;
  reg                 controlStream_s2mPipe_rData_firstRow;
  reg                 controlStream_s2mPipe_rData_lastRow;
  reg                 controlStream_s2mPipe_rData_finalResult;
  reg                 controlStream_s2mPipe_rData_mainCompare;
  reg                 controlStream_s2mPipe_rData_counterCompare;
  reg                 controlStream_s2mPipe_rData_horizontalCompare;
  reg                 controlStream_s2mPipe_rData_verticalCompare;
  reg        [7:0]    controlStream_s2mPipe_rData_mainDiff;
  reg        [7:0]    controlStream_s2mPipe_rData_counterDiff;
  reg        [7:0]    controlStream_s2mPipe_rData_horizontalDiff;
  reg        [7:0]    controlStream_s2mPipe_rData_verticalDiff;
  reg                 controlStream_s2mPipe_rData_isHorizontalMin;
  reg        [7:0]    controlStream_s2mPipe_rData_minDiff;
  reg        [1:0]    controlStream_s2mPipe_rData_currentPosition;
  reg        [1:0]    controlStream_s2mPipe_rData_nextPosition;
  reg                 controlStream_s2mPipe_rData_horizontalDirectionValid;
  reg                 controlStream_s2mPipe_rData_verticalDirectionValid;
  reg                 controlStream_s2mPipe_rData_mainDirectionValid;
  reg                 controlStream_s2mPipe_rData_counterDirectionValid;
  reg                 controlStream_s2mPipe_rData_inValidMinDiff;
  wire                when_Stream_l368_25;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_valid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_ready;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_frameStart;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_rowEnd;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_pipeValid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_firstRow;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_lastRow;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_finalResult;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainCompare;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterCompare;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_horizontalCompare;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_verticalCompare;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_horizontalDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_verticalDiff;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_isHorizontalMin;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_minDiff;
  wire       [1:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_currentPosition;
  wire       [1:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_nextPosition;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_horizontalDirectionValid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_verticalDirectionValid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDirectionValid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDirectionValid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_inValidMinDiff;
  reg                 controlStream_s2mPipe_m2sPipe_rValid;
  reg                 controlStream_s2mPipe_m2sPipe_rData_frameStart;
  reg                 controlStream_s2mPipe_m2sPipe_rData_rowEnd;
  reg                 controlStream_s2mPipe_m2sPipe_rData_pipeValid;
  reg                 controlStream_s2mPipe_m2sPipe_rData_firstRow;
  reg                 controlStream_s2mPipe_m2sPipe_rData_lastRow;
  reg                 controlStream_s2mPipe_m2sPipe_rData_finalResult;
  reg                 controlStream_s2mPipe_m2sPipe_rData_mainCompare;
  reg                 controlStream_s2mPipe_m2sPipe_rData_counterCompare;
  reg                 controlStream_s2mPipe_m2sPipe_rData_horizontalCompare;
  reg                 controlStream_s2mPipe_m2sPipe_rData_verticalCompare;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_rData_mainDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_rData_counterDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_rData_horizontalDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_rData_verticalDiff;
  reg                 controlStream_s2mPipe_m2sPipe_rData_isHorizontalMin;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_rData_minDiff;
  reg        [1:0]    controlStream_s2mPipe_m2sPipe_rData_currentPosition;
  reg        [1:0]    controlStream_s2mPipe_m2sPipe_rData_nextPosition;
  reg                 controlStream_s2mPipe_m2sPipe_rData_horizontalDirectionValid;
  reg                 controlStream_s2mPipe_m2sPipe_rData_verticalDirectionValid;
  reg                 controlStream_s2mPipe_m2sPipe_rData_mainDirectionValid;
  reg                 controlStream_s2mPipe_m2sPipe_rData_counterDirectionValid;
  reg                 controlStream_s2mPipe_m2sPipe_rData_inValidMinDiff;
  wire                when_Stream_l368_26;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_valid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_frameStart;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_rowEnd;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_pipeValid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_firstRow;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_lastRow;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_finalResult;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainCompare;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterCompare;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_horizontalCompare;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_verticalCompare;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_horizontalDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_verticalDiff;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_isHorizontalMin;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_minDiff;
  wire       [1:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_currentPosition;
  wire       [1:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_nextPosition;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_horizontalDirectionValid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_verticalDirectionValid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainDirectionValid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterDirectionValid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_inValidMinDiff;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_frameStart;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_rowEnd;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_pipeValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_firstRow;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_lastRow;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_finalResult;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainCompare;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterCompare;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_horizontalCompare;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_verticalCompare;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_horizontalDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_verticalDiff;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_isHorizontalMin;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_minDiff;
  reg        [1:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_currentPosition;
  reg        [1:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_nextPosition;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_horizontalDirectionValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_verticalDirectionValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainDirectionValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterDirectionValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_inValidMinDiff;
  wire                readStage_controlPipe_valid;
  wire                readStage_controlPipe_ready;
  wire                readStage_controlPipe_payload_frameStart;
  wire                readStage_controlPipe_payload_rowEnd;
  wire                readStage_controlPipe_payload_pipeValid;
  wire                readStage_controlPipe_payload_firstRow;
  wire                readStage_controlPipe_payload_lastRow;
  wire                readStage_controlPipe_payload_finalResult;
  wire                readStage_controlPipe_payload_mainCompare;
  wire                readStage_controlPipe_payload_counterCompare;
  wire                readStage_controlPipe_payload_horizontalCompare;
  wire                readStage_controlPipe_payload_verticalCompare;
  wire       [7:0]    readStage_controlPipe_payload_mainDiff;
  wire       [7:0]    readStage_controlPipe_payload_counterDiff;
  wire       [7:0]    readStage_controlPipe_payload_horizontalDiff;
  wire       [7:0]    readStage_controlPipe_payload_verticalDiff;
  wire                readStage_controlPipe_payload_isHorizontalMin;
  wire       [7:0]    readStage_controlPipe_payload_minDiff;
  wire       [1:0]    readStage_controlPipe_payload_currentPosition;
  wire       [1:0]    readStage_controlPipe_payload_nextPosition;
  wire                readStage_controlPipe_payload_horizontalDirectionValid;
  wire                readStage_controlPipe_payload_verticalDirectionValid;
  wire                readStage_controlPipe_payload_mainDirectionValid;
  wire                readStage_controlPipe_payload_counterDirectionValid;
  wire                readStage_controlPipe_payload_inValidMinDiff;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_frameStart;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_rowEnd;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_pipeValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_firstRow;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_lastRow;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_finalResult;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainCompare;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterCompare;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_horizontalCompare;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_verticalCompare;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_horizontalDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_verticalDiff;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_isHorizontalMin;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_minDiff;
  reg        [1:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_currentPosition;
  reg        [1:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_nextPosition;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_horizontalDirectionValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_verticalDirectionValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainDirectionValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterDirectionValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_inValidMinDiff;
  wire                when_Stream_l368_27;
  wire                readStage_mainOnePixelStream_s2mPipe_valid;
  reg                 readStage_mainOnePixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_mainOnePixelStream_s2mPipe_payload;
  reg                 readStage_mainOnePixelStream_rValid;
  reg        [7:0]    readStage_mainOnePixelStream_rData;
  wire                compareStage_mainOnePixelStream_valid;
  wire                compareStage_mainOnePixelStream_ready;
  wire       [7:0]    compareStage_mainOnePixelStream_payload;
  reg                 readStage_mainOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_mainOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_28;
  wire                readStage_counterOnePixelStream_s2mPipe_valid;
  reg                 readStage_counterOnePixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_counterOnePixelStream_s2mPipe_payload;
  reg                 readStage_counterOnePixelStream_rValid;
  reg        [7:0]    readStage_counterOnePixelStream_rData;
  wire                compareStage_counterOnePixelStream_valid;
  wire                compareStage_counterOnePixelStream_ready;
  wire       [7:0]    compareStage_counterOnePixelStream_payload;
  reg                 readStage_counterOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_counterOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_29;
  wire                readStage_mainTwoPixelStream_s2mPipe_valid;
  reg                 readStage_mainTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_mainTwoPixelStream_s2mPipe_payload;
  reg                 readStage_mainTwoPixelStream_rValid;
  reg        [7:0]    readStage_mainTwoPixelStream_rData;
  wire                compareStage_mainTwoPixelStream_valid;
  wire                compareStage_mainTwoPixelStream_ready;
  wire       [7:0]    compareStage_mainTwoPixelStream_payload;
  reg                 readStage_mainTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_mainTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_30;
  wire                readStage_counterTwoPixelStream_s2mPipe_valid;
  reg                 readStage_counterTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_counterTwoPixelStream_s2mPipe_payload;
  reg                 readStage_counterTwoPixelStream_rValid;
  reg        [7:0]    readStage_counterTwoPixelStream_rData;
  wire                compareStage_counterTwoPixelStream_valid;
  wire                compareStage_counterTwoPixelStream_ready;
  wire       [7:0]    compareStage_counterTwoPixelStream_payload;
  reg                 readStage_counterTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_counterTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_31;
  wire                readStage_mainThreePixelStream_s2mPipe_valid;
  reg                 readStage_mainThreePixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_mainThreePixelStream_s2mPipe_payload;
  reg                 readStage_mainThreePixelStream_rValid;
  reg        [7:0]    readStage_mainThreePixelStream_rData;
  wire                compareStage_mainThreePixelStream_valid;
  wire                compareStage_mainThreePixelStream_ready;
  wire       [7:0]    compareStage_mainThreePixelStream_payload;
  reg                 readStage_mainThreePixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_mainThreePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_32;
  wire                readStage_counterThreePixelStream_s2mPipe_valid;
  reg                 readStage_counterThreePixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_counterThreePixelStream_s2mPipe_payload;
  reg                 readStage_counterThreePixelStream_rValid;
  reg        [7:0]    readStage_counterThreePixelStream_rData;
  wire                compareStage_counterThreePixelStream_valid;
  wire                compareStage_counterThreePixelStream_ready;
  wire       [7:0]    compareStage_counterThreePixelStream_payload;
  reg                 readStage_counterThreePixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_counterThreePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_33;
  wire                readStage_mainOneValidStream_s2mPipe_valid;
  reg                 readStage_mainOneValidStream_s2mPipe_ready;
  wire                readStage_mainOneValidStream_s2mPipe_payload;
  reg                 readStage_mainOneValidStream_rValid;
  reg                 readStage_mainOneValidStream_rData;
  wire                compareStage_mainOneValidStream_valid;
  wire                compareStage_mainOneValidStream_ready;
  wire                compareStage_mainOneValidStream_payload;
  reg                 readStage_mainOneValidStream_s2mPipe_rValid;
  reg                 readStage_mainOneValidStream_s2mPipe_rData;
  wire                when_Stream_l368_34;
  wire                readStage_counterOneValidStream_s2mPipe_valid;
  reg                 readStage_counterOneValidStream_s2mPipe_ready;
  wire                readStage_counterOneValidStream_s2mPipe_payload;
  reg                 readStage_counterOneValidStream_rValid;
  reg                 readStage_counterOneValidStream_rData;
  wire                compareStage_counterOneValidStream_valid;
  wire                compareStage_counterOneValidStream_ready;
  wire                compareStage_counterOneValidStream_payload;
  reg                 readStage_counterOneValidStream_s2mPipe_rValid;
  reg                 readStage_counterOneValidStream_s2mPipe_rData;
  wire                when_Stream_l368_35;
  wire                readStage_mainTwoValidStream_s2mPipe_valid;
  reg                 readStage_mainTwoValidStream_s2mPipe_ready;
  wire                readStage_mainTwoValidStream_s2mPipe_payload;
  reg                 readStage_mainTwoValidStream_rValid;
  reg                 readStage_mainTwoValidStream_rData;
  wire                compareStage_mainTwoValidStream_valid;
  wire                compareStage_mainTwoValidStream_ready;
  wire                compareStage_mainTwoValidStream_payload;
  reg                 readStage_mainTwoValidStream_s2mPipe_rValid;
  reg                 readStage_mainTwoValidStream_s2mPipe_rData;
  wire                when_Stream_l368_36;
  wire                readStage_counterTwoValidStream_s2mPipe_valid;
  reg                 readStage_counterTwoValidStream_s2mPipe_ready;
  wire                readStage_counterTwoValidStream_s2mPipe_payload;
  reg                 readStage_counterTwoValidStream_rValid;
  reg                 readStage_counterTwoValidStream_rData;
  wire                compareStage_counterTwoValidStream_valid;
  wire                compareStage_counterTwoValidStream_ready;
  wire                compareStage_counterTwoValidStream_payload;
  reg                 readStage_counterTwoValidStream_s2mPipe_rValid;
  reg                 readStage_counterTwoValidStream_s2mPipe_rData;
  wire                when_Stream_l368_37;
  wire                readStage_mainThreeValidStream_s2mPipe_valid;
  reg                 readStage_mainThreeValidStream_s2mPipe_ready;
  wire                readStage_mainThreeValidStream_s2mPipe_payload;
  reg                 readStage_mainThreeValidStream_rValid;
  reg                 readStage_mainThreeValidStream_rData;
  wire                compareStage_mainThreeValidStream_valid;
  wire                compareStage_mainThreeValidStream_ready;
  wire                compareStage_mainThreeValidStream_payload;
  reg                 readStage_mainThreeValidStream_s2mPipe_rValid;
  reg                 readStage_mainThreeValidStream_s2mPipe_rData;
  wire                when_Stream_l368_38;
  wire                readStage_counterThreeValidStream_s2mPipe_valid;
  reg                 readStage_counterThreeValidStream_s2mPipe_ready;
  wire                readStage_counterThreeValidStream_s2mPipe_payload;
  reg                 readStage_counterThreeValidStream_rValid;
  reg                 readStage_counterThreeValidStream_rData;
  wire                compareStage_counterThreeValidStream_valid;
  wire                compareStage_counterThreeValidStream_ready;
  wire                compareStage_counterThreeValidStream_payload;
  reg                 readStage_counterThreeValidStream_s2mPipe_rValid;
  reg                 readStage_counterThreeValidStream_s2mPipe_rData;
  wire                when_Stream_l368_39;
  reg                 CICC1851_readStage_controlPipe_translated_payload_mainCompare;
  reg                 CICC1851_readStage_controlPipe_translated_payload_counterCompare;
  reg                 CICC1851_readStage_controlPipe_translated_payload_horizontalCompare;
  reg                 CICC1851_readStage_controlPipe_translated_payload_verticalCompare;
  reg                 CICC1851_readStage_controlPipe_translated_payload_horizontalDirectionValid;
  reg                 CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid;
  reg                 CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid;
  reg                 CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid;
  wire                when_SuperResolutionPart3_l342;
  wire                when_SuperResolutionPart3_l344;
  wire                when_SuperResolutionPart3_l345;
  wire                when_SuperResolutionPart3_l348;
  wire                when_SuperResolutionPart3_l351;
  wire                when_SuperResolutionPart3_l347;
  wire                when_SuperResolutionPart3_l356;
  wire                when_SuperResolutionPart3_l357;
  wire                when_SuperResolutionPart3_l365;
  wire                when_SuperResolutionPart3_l373;
  wire                when_SuperResolutionPart3_l378;
  wire                when_SuperResolutionPart3_l383;
  wire                when_SuperResolutionPart3_l391;
  wire                when_SuperResolutionPart3_l396;
  wire                when_SuperResolutionPart3_l401;
  wire                when_SuperResolutionPart3_l409;
  wire                when_SuperResolutionPart3_l377;
  wire                when_SuperResolutionPart3_l415;
  wire                when_SuperResolutionPart3_l416;
  wire                when_SuperResolutionPart3_l419;
  wire                when_SuperResolutionPart3_l422;
  wire                when_SuperResolutionPart3_l424;
  wire                when_SuperResolutionPart3_l432;
  wire                when_SuperResolutionPart3_l441;
  wire                when_SuperResolutionPart3_l449;
  wire                when_SuperResolutionPart3_l458;
  wire                when_SuperResolutionPart3_l460;
  wire                when_SuperResolutionPart3_l463;
  wire                when_SuperResolutionPart3_l465;
  wire                when_SuperResolutionPart3_l470;
  wire                when_SuperResolutionPart3_l477;
  wire                when_SuperResolutionPart3_l485;
  wire                when_SuperResolutionPart3_l487;
  wire                when_SuperResolutionPart3_l490;
  wire                when_SuperResolutionPart3_l492;
  wire                when_SuperResolutionPart3_l497;
  wire                when_SuperResolutionPart3_l500;
  wire                when_SuperResolutionPart3_l502;
  wire                when_SuperResolutionPart3_l504;
  wire                when_SuperResolutionPart3_l511;
  wire                when_SuperResolutionPart3_l519;
  wire                when_SuperResolutionPart3_l521;
  wire                when_SuperResolutionPart3_l524;
  wire                when_SuperResolutionPart3_l526;
  wire                when_SuperResolutionPart3_l531;
  wire                when_SuperResolutionPart3_l539;
  wire                when_SuperResolutionPart3_l547;
  wire                when_SuperResolutionPart3_l549;
  wire                when_SuperResolutionPart3_l552;
  wire                when_SuperResolutionPart3_l554;
  wire                when_SuperResolutionPart3_l559;
  wire                when_SuperResolutionPart3_l562;
  wire                when_SuperResolutionPart3_l564;
  wire                when_SuperResolutionPart3_l566;
  wire                when_SuperResolutionPart3_l573;
  wire                when_SuperResolutionPart3_l581;
  wire                when_SuperResolutionPart3_l583;
  wire                when_SuperResolutionPart3_l586;
  wire                when_SuperResolutionPart3_l588;
  wire                when_SuperResolutionPart3_l593;
  wire                when_SuperResolutionPart3_l601;
  wire                when_SuperResolutionPart3_l609;
  wire                when_SuperResolutionPart3_l611;
  wire                when_SuperResolutionPart3_l614;
  wire                when_SuperResolutionPart3_l616;
  wire                when_SuperResolutionPart3_l496;
  wire                readStage_controlPipe_translated_valid;
  wire                readStage_controlPipe_translated_ready;
  wire                readStage_controlPipe_translated_payload_frameStart;
  wire                readStage_controlPipe_translated_payload_rowEnd;
  wire                readStage_controlPipe_translated_payload_pipeValid;
  wire                readStage_controlPipe_translated_payload_firstRow;
  wire                readStage_controlPipe_translated_payload_lastRow;
  wire                readStage_controlPipe_translated_payload_finalResult;
  wire                readStage_controlPipe_translated_payload_mainCompare;
  wire                readStage_controlPipe_translated_payload_counterCompare;
  wire                readStage_controlPipe_translated_payload_horizontalCompare;
  wire                readStage_controlPipe_translated_payload_verticalCompare;
  wire       [7:0]    readStage_controlPipe_translated_payload_mainDiff;
  wire       [7:0]    readStage_controlPipe_translated_payload_counterDiff;
  wire       [7:0]    readStage_controlPipe_translated_payload_horizontalDiff;
  wire       [7:0]    readStage_controlPipe_translated_payload_verticalDiff;
  wire                readStage_controlPipe_translated_payload_isHorizontalMin;
  wire       [7:0]    readStage_controlPipe_translated_payload_minDiff;
  wire       [1:0]    readStage_controlPipe_translated_payload_currentPosition;
  wire       [1:0]    readStage_controlPipe_translated_payload_nextPosition;
  wire                readStage_controlPipe_translated_payload_horizontalDirectionValid;
  wire                readStage_controlPipe_translated_payload_verticalDirectionValid;
  wire                readStage_controlPipe_translated_payload_mainDirectionValid;
  wire                readStage_controlPipe_translated_payload_counterDirectionValid;
  wire                readStage_controlPipe_translated_payload_inValidMinDiff;
  wire                readStage_controlPipe_translated_s2mPipe_valid;
  reg                 readStage_controlPipe_translated_s2mPipe_ready;
  wire                readStage_controlPipe_translated_s2mPipe_payload_frameStart;
  wire                readStage_controlPipe_translated_s2mPipe_payload_rowEnd;
  wire                readStage_controlPipe_translated_s2mPipe_payload_pipeValid;
  wire                readStage_controlPipe_translated_s2mPipe_payload_firstRow;
  wire                readStage_controlPipe_translated_s2mPipe_payload_lastRow;
  wire                readStage_controlPipe_translated_s2mPipe_payload_finalResult;
  wire                readStage_controlPipe_translated_s2mPipe_payload_mainCompare;
  wire                readStage_controlPipe_translated_s2mPipe_payload_counterCompare;
  wire                readStage_controlPipe_translated_s2mPipe_payload_horizontalCompare;
  wire                readStage_controlPipe_translated_s2mPipe_payload_verticalCompare;
  wire       [7:0]    readStage_controlPipe_translated_s2mPipe_payload_mainDiff;
  wire       [7:0]    readStage_controlPipe_translated_s2mPipe_payload_counterDiff;
  wire       [7:0]    readStage_controlPipe_translated_s2mPipe_payload_horizontalDiff;
  wire       [7:0]    readStage_controlPipe_translated_s2mPipe_payload_verticalDiff;
  wire                readStage_controlPipe_translated_s2mPipe_payload_isHorizontalMin;
  wire       [7:0]    readStage_controlPipe_translated_s2mPipe_payload_minDiff;
  wire       [1:0]    readStage_controlPipe_translated_s2mPipe_payload_currentPosition;
  wire       [1:0]    readStage_controlPipe_translated_s2mPipe_payload_nextPosition;
  wire                readStage_controlPipe_translated_s2mPipe_payload_horizontalDirectionValid;
  wire                readStage_controlPipe_translated_s2mPipe_payload_verticalDirectionValid;
  wire                readStage_controlPipe_translated_s2mPipe_payload_mainDirectionValid;
  wire                readStage_controlPipe_translated_s2mPipe_payload_counterDirectionValid;
  wire                readStage_controlPipe_translated_s2mPipe_payload_inValidMinDiff;
  reg                 readStage_controlPipe_translated_rValid;
  reg                 readStage_controlPipe_translated_rData_frameStart;
  reg                 readStage_controlPipe_translated_rData_rowEnd;
  reg                 readStage_controlPipe_translated_rData_pipeValid;
  reg                 readStage_controlPipe_translated_rData_firstRow;
  reg                 readStage_controlPipe_translated_rData_lastRow;
  reg                 readStage_controlPipe_translated_rData_finalResult;
  reg                 readStage_controlPipe_translated_rData_mainCompare;
  reg                 readStage_controlPipe_translated_rData_counterCompare;
  reg                 readStage_controlPipe_translated_rData_horizontalCompare;
  reg                 readStage_controlPipe_translated_rData_verticalCompare;
  reg        [7:0]    readStage_controlPipe_translated_rData_mainDiff;
  reg        [7:0]    readStage_controlPipe_translated_rData_counterDiff;
  reg        [7:0]    readStage_controlPipe_translated_rData_horizontalDiff;
  reg        [7:0]    readStage_controlPipe_translated_rData_verticalDiff;
  reg                 readStage_controlPipe_translated_rData_isHorizontalMin;
  reg        [7:0]    readStage_controlPipe_translated_rData_minDiff;
  reg        [1:0]    readStage_controlPipe_translated_rData_currentPosition;
  reg        [1:0]    readStage_controlPipe_translated_rData_nextPosition;
  reg                 readStage_controlPipe_translated_rData_horizontalDirectionValid;
  reg                 readStage_controlPipe_translated_rData_verticalDirectionValid;
  reg                 readStage_controlPipe_translated_rData_mainDirectionValid;
  reg                 readStage_controlPipe_translated_rData_counterDirectionValid;
  reg                 readStage_controlPipe_translated_rData_inValidMinDiff;
  wire                compareStage_controlPipe_valid;
  wire                compareStage_controlPipe_ready;
  wire                compareStage_controlPipe_payload_frameStart;
  wire                compareStage_controlPipe_payload_rowEnd;
  wire                compareStage_controlPipe_payload_pipeValid;
  wire                compareStage_controlPipe_payload_firstRow;
  wire                compareStage_controlPipe_payload_lastRow;
  wire                compareStage_controlPipe_payload_finalResult;
  wire                compareStage_controlPipe_payload_mainCompare;
  wire                compareStage_controlPipe_payload_counterCompare;
  wire                compareStage_controlPipe_payload_horizontalCompare;
  wire                compareStage_controlPipe_payload_verticalCompare;
  wire       [7:0]    compareStage_controlPipe_payload_mainDiff;
  wire       [7:0]    compareStage_controlPipe_payload_counterDiff;
  wire       [7:0]    compareStage_controlPipe_payload_horizontalDiff;
  wire       [7:0]    compareStage_controlPipe_payload_verticalDiff;
  wire                compareStage_controlPipe_payload_isHorizontalMin;
  wire       [7:0]    compareStage_controlPipe_payload_minDiff;
  wire       [1:0]    compareStage_controlPipe_payload_currentPosition;
  wire       [1:0]    compareStage_controlPipe_payload_nextPosition;
  wire                compareStage_controlPipe_payload_horizontalDirectionValid;
  wire                compareStage_controlPipe_payload_verticalDirectionValid;
  wire                compareStage_controlPipe_payload_mainDirectionValid;
  wire                compareStage_controlPipe_payload_counterDirectionValid;
  wire                compareStage_controlPipe_payload_inValidMinDiff;
  reg                 readStage_controlPipe_translated_s2mPipe_rValid;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_frameStart;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_rowEnd;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_pipeValid;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_firstRow;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_lastRow;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_finalResult;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_mainCompare;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_counterCompare;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_horizontalCompare;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_verticalCompare;
  reg        [7:0]    readStage_controlPipe_translated_s2mPipe_rData_mainDiff;
  reg        [7:0]    readStage_controlPipe_translated_s2mPipe_rData_counterDiff;
  reg        [7:0]    readStage_controlPipe_translated_s2mPipe_rData_horizontalDiff;
  reg        [7:0]    readStage_controlPipe_translated_s2mPipe_rData_verticalDiff;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_isHorizontalMin;
  reg        [7:0]    readStage_controlPipe_translated_s2mPipe_rData_minDiff;
  reg        [1:0]    readStage_controlPipe_translated_s2mPipe_rData_currentPosition;
  reg        [1:0]    readStage_controlPipe_translated_s2mPipe_rData_nextPosition;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_horizontalDirectionValid;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_verticalDirectionValid;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_mainDirectionValid;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_counterDirectionValid;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_inValidMinDiff;
  wire                when_Stream_l368_40;
  wire                compareStage_mainOnePixelStream_s2mPipe_valid;
  reg                 compareStage_mainOnePixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_mainOnePixelStream_s2mPipe_payload;
  reg                 compareStage_mainOnePixelStream_rValid;
  reg        [7:0]    compareStage_mainOnePixelStream_rData;
  wire                diffStage_mainOnePixelStream_valid;
  wire                diffStage_mainOnePixelStream_ready;
  wire       [7:0]    diffStage_mainOnePixelStream_payload;
  reg                 compareStage_mainOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_mainOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_41;
  wire                compareStage_counterOnePixelStream_s2mPipe_valid;
  reg                 compareStage_counterOnePixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_counterOnePixelStream_s2mPipe_payload;
  reg                 compareStage_counterOnePixelStream_rValid;
  reg        [7:0]    compareStage_counterOnePixelStream_rData;
  wire                diffStage_counterOnePixelStream_valid;
  wire                diffStage_counterOnePixelStream_ready;
  wire       [7:0]    diffStage_counterOnePixelStream_payload;
  reg                 compareStage_counterOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_counterOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_42;
  wire                compareStage_mainTwoPixelStream_s2mPipe_valid;
  reg                 compareStage_mainTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_mainTwoPixelStream_s2mPipe_payload;
  reg                 compareStage_mainTwoPixelStream_rValid;
  reg        [7:0]    compareStage_mainTwoPixelStream_rData;
  wire                diffStage_mainTwoPixelStream_valid;
  wire                diffStage_mainTwoPixelStream_ready;
  wire       [7:0]    diffStage_mainTwoPixelStream_payload;
  reg                 compareStage_mainTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_mainTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_43;
  wire                compareStage_counterTwoPixelStream_s2mPipe_valid;
  reg                 compareStage_counterTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_counterTwoPixelStream_s2mPipe_payload;
  reg                 compareStage_counterTwoPixelStream_rValid;
  reg        [7:0]    compareStage_counterTwoPixelStream_rData;
  wire                diffStage_counterTwoPixelStream_valid;
  wire                diffStage_counterTwoPixelStream_ready;
  wire       [7:0]    diffStage_counterTwoPixelStream_payload;
  reg                 compareStage_counterTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_counterTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_44;
  wire                compareStage_mainThreePixelStream_s2mPipe_valid;
  reg                 compareStage_mainThreePixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_mainThreePixelStream_s2mPipe_payload;
  reg                 compareStage_mainThreePixelStream_rValid;
  reg        [7:0]    compareStage_mainThreePixelStream_rData;
  wire                diffStage_mainThreePixelStream_valid;
  wire                diffStage_mainThreePixelStream_ready;
  wire       [7:0]    diffStage_mainThreePixelStream_payload;
  reg                 compareStage_mainThreePixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_mainThreePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_45;
  wire                compareStage_counterThreePixelStream_s2mPipe_valid;
  reg                 compareStage_counterThreePixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_counterThreePixelStream_s2mPipe_payload;
  reg                 compareStage_counterThreePixelStream_rValid;
  reg        [7:0]    compareStage_counterThreePixelStream_rData;
  wire                diffStage_counterThreePixelStream_valid;
  wire                diffStage_counterThreePixelStream_ready;
  wire       [7:0]    diffStage_counterThreePixelStream_payload;
  reg                 compareStage_counterThreePixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_counterThreePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_46;
  wire                compareStage_mainOneValidStream_s2mPipe_valid;
  reg                 compareStage_mainOneValidStream_s2mPipe_ready;
  wire                compareStage_mainOneValidStream_s2mPipe_payload;
  reg                 compareStage_mainOneValidStream_rValid;
  reg                 compareStage_mainOneValidStream_rData;
  wire                diffStage_mainOneValidStream_valid;
  wire                diffStage_mainOneValidStream_ready;
  wire                diffStage_mainOneValidStream_payload;
  reg                 compareStage_mainOneValidStream_s2mPipe_rValid;
  reg                 compareStage_mainOneValidStream_s2mPipe_rData;
  wire                when_Stream_l368_47;
  wire                compareStage_counterOneValidStream_s2mPipe_valid;
  reg                 compareStage_counterOneValidStream_s2mPipe_ready;
  wire                compareStage_counterOneValidStream_s2mPipe_payload;
  reg                 compareStage_counterOneValidStream_rValid;
  reg                 compareStage_counterOneValidStream_rData;
  wire                diffStage_counterOneValidStream_valid;
  wire                diffStage_counterOneValidStream_ready;
  wire                diffStage_counterOneValidStream_payload;
  reg                 compareStage_counterOneValidStream_s2mPipe_rValid;
  reg                 compareStage_counterOneValidStream_s2mPipe_rData;
  wire                when_Stream_l368_48;
  wire                compareStage_mainTwoValidStream_s2mPipe_valid;
  reg                 compareStage_mainTwoValidStream_s2mPipe_ready;
  wire                compareStage_mainTwoValidStream_s2mPipe_payload;
  reg                 compareStage_mainTwoValidStream_rValid;
  reg                 compareStage_mainTwoValidStream_rData;
  wire                diffStage_mainTwoValidStream_valid;
  wire                diffStage_mainTwoValidStream_ready;
  wire                diffStage_mainTwoValidStream_payload;
  reg                 compareStage_mainTwoValidStream_s2mPipe_rValid;
  reg                 compareStage_mainTwoValidStream_s2mPipe_rData;
  wire                when_Stream_l368_49;
  wire                compareStage_counterTwoValidStream_s2mPipe_valid;
  reg                 compareStage_counterTwoValidStream_s2mPipe_ready;
  wire                compareStage_counterTwoValidStream_s2mPipe_payload;
  reg                 compareStage_counterTwoValidStream_rValid;
  reg                 compareStage_counterTwoValidStream_rData;
  wire                diffStage_counterTwoValidStream_valid;
  wire                diffStage_counterTwoValidStream_ready;
  wire                diffStage_counterTwoValidStream_payload;
  reg                 compareStage_counterTwoValidStream_s2mPipe_rValid;
  reg                 compareStage_counterTwoValidStream_s2mPipe_rData;
  wire                when_Stream_l368_50;
  wire                compareStage_mainThreeValidStream_s2mPipe_valid;
  reg                 compareStage_mainThreeValidStream_s2mPipe_ready;
  wire                compareStage_mainThreeValidStream_s2mPipe_payload;
  reg                 compareStage_mainThreeValidStream_rValid;
  reg                 compareStage_mainThreeValidStream_rData;
  wire                diffStage_mainThreeValidStream_valid;
  wire                diffStage_mainThreeValidStream_ready;
  wire                diffStage_mainThreeValidStream_payload;
  reg                 compareStage_mainThreeValidStream_s2mPipe_rValid;
  reg                 compareStage_mainThreeValidStream_s2mPipe_rData;
  wire                when_Stream_l368_51;
  wire                compareStage_counterThreeValidStream_s2mPipe_valid;
  reg                 compareStage_counterThreeValidStream_s2mPipe_ready;
  wire                compareStage_counterThreeValidStream_s2mPipe_payload;
  reg                 compareStage_counterThreeValidStream_rValid;
  reg                 compareStage_counterThreeValidStream_rData;
  wire                diffStage_counterThreeValidStream_valid;
  wire                diffStage_counterThreeValidStream_ready;
  wire                diffStage_counterThreeValidStream_payload;
  reg                 compareStage_counterThreeValidStream_s2mPipe_rValid;
  reg                 compareStage_counterThreeValidStream_s2mPipe_rData;
  wire                when_Stream_l368_52;
  reg        [7:0]    CICC1851_compareStage_controlPipe_translated_payload_mainDiff;
  reg        [7:0]    CICC1851_compareStage_controlPipe_translated_payload_counterDiff;
  reg        [7:0]    CICC1851_compareStage_controlPipe_translated_payload_horizontalDiff;
  reg        [7:0]    CICC1851_compareStage_controlPipe_translated_payload_verticalDiff;
  reg                 CICC1851_compareStage_controlPipe_translated_payload_inValidMinDiff;
  wire                when_SuperResolutionPart3_l647;
  wire                when_SuperResolutionPart3_l649;
  wire                when_SuperResolutionPart3_l652;
  wire                when_SuperResolutionPart3_l661;
  wire                when_SuperResolutionPart3_l664;
  wire                when_SuperResolutionPart3_l697;
  wire                when_SuperResolutionPart3_l725;
  wire                when_SuperResolutionPart3_l694;
  wire                when_SuperResolutionPart3_l753;
  wire                compareStage_controlPipe_translated_valid;
  wire                compareStage_controlPipe_translated_ready;
  wire                compareStage_controlPipe_translated_payload_frameStart;
  wire                compareStage_controlPipe_translated_payload_rowEnd;
  wire                compareStage_controlPipe_translated_payload_pipeValid;
  wire                compareStage_controlPipe_translated_payload_firstRow;
  wire                compareStage_controlPipe_translated_payload_lastRow;
  wire                compareStage_controlPipe_translated_payload_finalResult;
  wire                compareStage_controlPipe_translated_payload_mainCompare;
  wire                compareStage_controlPipe_translated_payload_counterCompare;
  wire                compareStage_controlPipe_translated_payload_horizontalCompare;
  wire                compareStage_controlPipe_translated_payload_verticalCompare;
  wire       [7:0]    compareStage_controlPipe_translated_payload_mainDiff;
  wire       [7:0]    compareStage_controlPipe_translated_payload_counterDiff;
  wire       [7:0]    compareStage_controlPipe_translated_payload_horizontalDiff;
  wire       [7:0]    compareStage_controlPipe_translated_payload_verticalDiff;
  wire                compareStage_controlPipe_translated_payload_isHorizontalMin;
  wire       [7:0]    compareStage_controlPipe_translated_payload_minDiff;
  wire       [1:0]    compareStage_controlPipe_translated_payload_currentPosition;
  wire       [1:0]    compareStage_controlPipe_translated_payload_nextPosition;
  wire                compareStage_controlPipe_translated_payload_horizontalDirectionValid;
  wire                compareStage_controlPipe_translated_payload_verticalDirectionValid;
  wire                compareStage_controlPipe_translated_payload_mainDirectionValid;
  wire                compareStage_controlPipe_translated_payload_counterDirectionValid;
  wire                compareStage_controlPipe_translated_payload_inValidMinDiff;
  wire                compareStage_controlPipe_translated_s2mPipe_valid;
  reg                 compareStage_controlPipe_translated_s2mPipe_ready;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_frameStart;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_rowEnd;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_pipeValid;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_firstRow;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_lastRow;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_finalResult;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_mainCompare;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_counterCompare;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_horizontalCompare;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_verticalCompare;
  wire       [7:0]    compareStage_controlPipe_translated_s2mPipe_payload_mainDiff;
  wire       [7:0]    compareStage_controlPipe_translated_s2mPipe_payload_counterDiff;
  wire       [7:0]    compareStage_controlPipe_translated_s2mPipe_payload_horizontalDiff;
  wire       [7:0]    compareStage_controlPipe_translated_s2mPipe_payload_verticalDiff;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_isHorizontalMin;
  wire       [7:0]    compareStage_controlPipe_translated_s2mPipe_payload_minDiff;
  wire       [1:0]    compareStage_controlPipe_translated_s2mPipe_payload_currentPosition;
  wire       [1:0]    compareStage_controlPipe_translated_s2mPipe_payload_nextPosition;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_horizontalDirectionValid;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_verticalDirectionValid;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_mainDirectionValid;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_counterDirectionValid;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_inValidMinDiff;
  reg                 compareStage_controlPipe_translated_rValid;
  reg                 compareStage_controlPipe_translated_rData_frameStart;
  reg                 compareStage_controlPipe_translated_rData_rowEnd;
  reg                 compareStage_controlPipe_translated_rData_pipeValid;
  reg                 compareStage_controlPipe_translated_rData_firstRow;
  reg                 compareStage_controlPipe_translated_rData_lastRow;
  reg                 compareStage_controlPipe_translated_rData_finalResult;
  reg                 compareStage_controlPipe_translated_rData_mainCompare;
  reg                 compareStage_controlPipe_translated_rData_counterCompare;
  reg                 compareStage_controlPipe_translated_rData_horizontalCompare;
  reg                 compareStage_controlPipe_translated_rData_verticalCompare;
  reg        [7:0]    compareStage_controlPipe_translated_rData_mainDiff;
  reg        [7:0]    compareStage_controlPipe_translated_rData_counterDiff;
  reg        [7:0]    compareStage_controlPipe_translated_rData_horizontalDiff;
  reg        [7:0]    compareStage_controlPipe_translated_rData_verticalDiff;
  reg                 compareStage_controlPipe_translated_rData_isHorizontalMin;
  reg        [7:0]    compareStage_controlPipe_translated_rData_minDiff;
  reg        [1:0]    compareStage_controlPipe_translated_rData_currentPosition;
  reg        [1:0]    compareStage_controlPipe_translated_rData_nextPosition;
  reg                 compareStage_controlPipe_translated_rData_horizontalDirectionValid;
  reg                 compareStage_controlPipe_translated_rData_verticalDirectionValid;
  reg                 compareStage_controlPipe_translated_rData_mainDirectionValid;
  reg                 compareStage_controlPipe_translated_rData_counterDirectionValid;
  reg                 compareStage_controlPipe_translated_rData_inValidMinDiff;
  wire                diffStage_controlPipe_valid;
  wire                diffStage_controlPipe_ready;
  wire                diffStage_controlPipe_payload_frameStart;
  wire                diffStage_controlPipe_payload_rowEnd;
  wire                diffStage_controlPipe_payload_pipeValid;
  wire                diffStage_controlPipe_payload_firstRow;
  wire                diffStage_controlPipe_payload_lastRow;
  wire                diffStage_controlPipe_payload_finalResult;
  wire                diffStage_controlPipe_payload_mainCompare;
  wire                diffStage_controlPipe_payload_counterCompare;
  wire                diffStage_controlPipe_payload_horizontalCompare;
  wire                diffStage_controlPipe_payload_verticalCompare;
  wire       [7:0]    diffStage_controlPipe_payload_mainDiff;
  wire       [7:0]    diffStage_controlPipe_payload_counterDiff;
  wire       [7:0]    diffStage_controlPipe_payload_horizontalDiff;
  wire       [7:0]    diffStage_controlPipe_payload_verticalDiff;
  wire                diffStage_controlPipe_payload_isHorizontalMin;
  wire       [7:0]    diffStage_controlPipe_payload_minDiff;
  wire       [1:0]    diffStage_controlPipe_payload_currentPosition;
  wire       [1:0]    diffStage_controlPipe_payload_nextPosition;
  wire                diffStage_controlPipe_payload_horizontalDirectionValid;
  wire                diffStage_controlPipe_payload_verticalDirectionValid;
  wire                diffStage_controlPipe_payload_mainDirectionValid;
  wire                diffStage_controlPipe_payload_counterDirectionValid;
  wire                diffStage_controlPipe_payload_inValidMinDiff;
  reg                 compareStage_controlPipe_translated_s2mPipe_rValid;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_frameStart;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_rowEnd;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_pipeValid;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_firstRow;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_lastRow;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_finalResult;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_mainCompare;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_counterCompare;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_horizontalCompare;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_verticalCompare;
  reg        [7:0]    compareStage_controlPipe_translated_s2mPipe_rData_mainDiff;
  reg        [7:0]    compareStage_controlPipe_translated_s2mPipe_rData_counterDiff;
  reg        [7:0]    compareStage_controlPipe_translated_s2mPipe_rData_horizontalDiff;
  reg        [7:0]    compareStage_controlPipe_translated_s2mPipe_rData_verticalDiff;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_isHorizontalMin;
  reg        [7:0]    compareStage_controlPipe_translated_s2mPipe_rData_minDiff;
  reg        [1:0]    compareStage_controlPipe_translated_s2mPipe_rData_currentPosition;
  reg        [1:0]    compareStage_controlPipe_translated_s2mPipe_rData_nextPosition;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_horizontalDirectionValid;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_verticalDirectionValid;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_mainDirectionValid;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_counterDirectionValid;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_inValidMinDiff;
  wire                when_Stream_l368_53;
  wire                diffStage_mainOnePixelStream_s2mPipe_valid;
  reg                 diffStage_mainOnePixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_mainOnePixelStream_s2mPipe_payload;
  reg                 diffStage_mainOnePixelStream_rValid;
  reg        [7:0]    diffStage_mainOnePixelStream_rData;
  wire                resultStage_mainOnePixelStream_valid;
  wire                resultStage_mainOnePixelStream_ready;
  wire       [7:0]    resultStage_mainOnePixelStream_payload;
  reg                 diffStage_mainOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_mainOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_54;
  wire                diffStage_counterOnePixelStream_s2mPipe_valid;
  reg                 diffStage_counterOnePixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_counterOnePixelStream_s2mPipe_payload;
  reg                 diffStage_counterOnePixelStream_rValid;
  reg        [7:0]    diffStage_counterOnePixelStream_rData;
  wire                resultStage_counterOnePixelStream_valid;
  wire                resultStage_counterOnePixelStream_ready;
  wire       [7:0]    resultStage_counterOnePixelStream_payload;
  reg                 diffStage_counterOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_counterOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_55;
  wire                diffStage_mainTwoPixelStream_s2mPipe_valid;
  reg                 diffStage_mainTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_mainTwoPixelStream_s2mPipe_payload;
  reg                 diffStage_mainTwoPixelStream_rValid;
  reg        [7:0]    diffStage_mainTwoPixelStream_rData;
  wire                resultStage_mainTwoPixelStream_valid;
  wire                resultStage_mainTwoPixelStream_ready;
  wire       [7:0]    resultStage_mainTwoPixelStream_payload;
  reg                 diffStage_mainTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_mainTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_56;
  wire                diffStage_counterTwoPixelStream_s2mPipe_valid;
  reg                 diffStage_counterTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_counterTwoPixelStream_s2mPipe_payload;
  reg                 diffStage_counterTwoPixelStream_rValid;
  reg        [7:0]    diffStage_counterTwoPixelStream_rData;
  wire                resultStage_counterTwoPixelStream_valid;
  wire                resultStage_counterTwoPixelStream_ready;
  wire       [7:0]    resultStage_counterTwoPixelStream_payload;
  reg                 diffStage_counterTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_counterTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_57;
  wire                diffStage_mainThreePixelStream_s2mPipe_valid;
  reg                 diffStage_mainThreePixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_mainThreePixelStream_s2mPipe_payload;
  reg                 diffStage_mainThreePixelStream_rValid;
  reg        [7:0]    diffStage_mainThreePixelStream_rData;
  wire                resultStage_mainThreePixelStream_valid;
  wire                resultStage_mainThreePixelStream_ready;
  wire       [7:0]    resultStage_mainThreePixelStream_payload;
  reg                 diffStage_mainThreePixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_mainThreePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_58;
  wire                diffStage_counterThreePixelStream_s2mPipe_valid;
  reg                 diffStage_counterThreePixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_counterThreePixelStream_s2mPipe_payload;
  reg                 diffStage_counterThreePixelStream_rValid;
  reg        [7:0]    diffStage_counterThreePixelStream_rData;
  wire                resultStage_counterThreePixelStream_valid;
  wire                resultStage_counterThreePixelStream_ready;
  wire       [7:0]    resultStage_counterThreePixelStream_payload;
  reg                 diffStage_counterThreePixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_counterThreePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_59;
  wire                diffStage_mainOneValidStream_s2mPipe_valid;
  reg                 diffStage_mainOneValidStream_s2mPipe_ready;
  wire                diffStage_mainOneValidStream_s2mPipe_payload;
  reg                 diffStage_mainOneValidStream_rValid;
  reg                 diffStage_mainOneValidStream_rData;
  wire                resultStage_mainOneValidStream_valid;
  wire                resultStage_mainOneValidStream_ready;
  wire                resultStage_mainOneValidStream_payload;
  reg                 diffStage_mainOneValidStream_s2mPipe_rValid;
  reg                 diffStage_mainOneValidStream_s2mPipe_rData;
  wire                when_Stream_l368_60;
  wire                diffStage_counterOneValidStream_s2mPipe_valid;
  reg                 diffStage_counterOneValidStream_s2mPipe_ready;
  wire                diffStage_counterOneValidStream_s2mPipe_payload;
  reg                 diffStage_counterOneValidStream_rValid;
  reg                 diffStage_counterOneValidStream_rData;
  wire                resultStage_counterOneValidStream_valid;
  wire                resultStage_counterOneValidStream_ready;
  wire                resultStage_counterOneValidStream_payload;
  reg                 diffStage_counterOneValidStream_s2mPipe_rValid;
  reg                 diffStage_counterOneValidStream_s2mPipe_rData;
  wire                when_Stream_l368_61;
  wire                diffStage_mainTwoValidStream_s2mPipe_valid;
  reg                 diffStage_mainTwoValidStream_s2mPipe_ready;
  wire                diffStage_mainTwoValidStream_s2mPipe_payload;
  reg                 diffStage_mainTwoValidStream_rValid;
  reg                 diffStage_mainTwoValidStream_rData;
  wire                resultStage_mainTwoValidStream_valid;
  wire                resultStage_mainTwoValidStream_ready;
  wire                resultStage_mainTwoValidStream_payload;
  reg                 diffStage_mainTwoValidStream_s2mPipe_rValid;
  reg                 diffStage_mainTwoValidStream_s2mPipe_rData;
  wire                when_Stream_l368_62;
  wire                diffStage_counterTwoValidStream_s2mPipe_valid;
  reg                 diffStage_counterTwoValidStream_s2mPipe_ready;
  wire                diffStage_counterTwoValidStream_s2mPipe_payload;
  reg                 diffStage_counterTwoValidStream_rValid;
  reg                 diffStage_counterTwoValidStream_rData;
  wire                resultStage_counterTwoValidStream_valid;
  wire                resultStage_counterTwoValidStream_ready;
  wire                resultStage_counterTwoValidStream_payload;
  reg                 diffStage_counterTwoValidStream_s2mPipe_rValid;
  reg                 diffStage_counterTwoValidStream_s2mPipe_rData;
  wire                when_Stream_l368_63;
  wire                diffStage_mainThreeValidStream_s2mPipe_valid;
  reg                 diffStage_mainThreeValidStream_s2mPipe_ready;
  wire                diffStage_mainThreeValidStream_s2mPipe_payload;
  reg                 diffStage_mainThreeValidStream_rValid;
  reg                 diffStage_mainThreeValidStream_rData;
  wire                resultStage_mainThreeValidStream_valid;
  wire                resultStage_mainThreeValidStream_ready;
  wire                resultStage_mainThreeValidStream_payload;
  reg                 diffStage_mainThreeValidStream_s2mPipe_rValid;
  reg                 diffStage_mainThreeValidStream_s2mPipe_rData;
  wire                when_Stream_l368_64;
  wire                diffStage_counterThreeValidStream_s2mPipe_valid;
  reg                 diffStage_counterThreeValidStream_s2mPipe_ready;
  wire                diffStage_counterThreeValidStream_s2mPipe_payload;
  reg                 diffStage_counterThreeValidStream_rValid;
  reg                 diffStage_counterThreeValidStream_rData;
  wire                resultStage_counterThreeValidStream_valid;
  wire                resultStage_counterThreeValidStream_ready;
  wire                resultStage_counterThreeValidStream_payload;
  reg                 diffStage_counterThreeValidStream_s2mPipe_rValid;
  reg                 diffStage_counterThreeValidStream_s2mPipe_rData;
  wire                when_Stream_l368_65;
  reg                 CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin;
  reg        [7:0]    CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff;
  wire                when_SuperResolutionPart3_l783;
  wire                when_SuperResolutionPart3_l784;
  wire                when_SuperResolutionPart3_l785;
  wire                when_SuperResolutionPart3_l788;
  wire                when_SuperResolutionPart3_l796;
  wire                when_SuperResolutionPart3_l804;
  wire                when_SuperResolutionPart3_l812;
  wire                when_SuperResolutionPart3_l795;
  wire                when_SuperResolutionPart3_l803;
  wire                when_SuperResolutionPart3_l811;
  wire                when_SuperResolutionPart3_l819;
  wire                when_SuperResolutionPart3_l822;
  wire                when_SuperResolutionPart3_l825;
  wire                resultStage_controlPipeBeforePipe_valid;
  wire                resultStage_controlPipeBeforePipe_ready;
  wire                resultStage_controlPipeBeforePipe_payload_frameStart;
  wire                resultStage_controlPipeBeforePipe_payload_rowEnd;
  wire                resultStage_controlPipeBeforePipe_payload_pipeValid;
  wire                resultStage_controlPipeBeforePipe_payload_firstRow;
  wire                resultStage_controlPipeBeforePipe_payload_lastRow;
  wire                resultStage_controlPipeBeforePipe_payload_finalResult;
  wire                resultStage_controlPipeBeforePipe_payload_mainCompare;
  wire                resultStage_controlPipeBeforePipe_payload_counterCompare;
  wire                resultStage_controlPipeBeforePipe_payload_horizontalCompare;
  wire                resultStage_controlPipeBeforePipe_payload_verticalCompare;
  wire       [7:0]    resultStage_controlPipeBeforePipe_payload_mainDiff;
  wire       [7:0]    resultStage_controlPipeBeforePipe_payload_counterDiff;
  wire       [7:0]    resultStage_controlPipeBeforePipe_payload_horizontalDiff;
  wire       [7:0]    resultStage_controlPipeBeforePipe_payload_verticalDiff;
  wire                resultStage_controlPipeBeforePipe_payload_isHorizontalMin;
  wire       [7:0]    resultStage_controlPipeBeforePipe_payload_minDiff;
  wire       [1:0]    resultStage_controlPipeBeforePipe_payload_currentPosition;
  wire       [1:0]    resultStage_controlPipeBeforePipe_payload_nextPosition;
  wire                resultStage_controlPipeBeforePipe_payload_horizontalDirectionValid;
  wire                resultStage_controlPipeBeforePipe_payload_verticalDirectionValid;
  wire                resultStage_controlPipeBeforePipe_payload_mainDirectionValid;
  wire                resultStage_controlPipeBeforePipe_payload_counterDirectionValid;
  wire                resultStage_controlPipeBeforePipe_payload_inValidMinDiff;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_valid;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_ready;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_frameStart;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_rowEnd;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_pipeValid;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_firstRow;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_lastRow;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_finalResult;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_mainCompare;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_counterCompare;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_horizontalCompare;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_verticalCompare;
  wire       [7:0]    resultStage_controlPipeBeforePipe_s2mPipe_payload_mainDiff;
  wire       [7:0]    resultStage_controlPipeBeforePipe_s2mPipe_payload_counterDiff;
  wire       [7:0]    resultStage_controlPipeBeforePipe_s2mPipe_payload_horizontalDiff;
  wire       [7:0]    resultStage_controlPipeBeforePipe_s2mPipe_payload_verticalDiff;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_isHorizontalMin;
  wire       [7:0]    resultStage_controlPipeBeforePipe_s2mPipe_payload_minDiff;
  wire       [1:0]    resultStage_controlPipeBeforePipe_s2mPipe_payload_currentPosition;
  wire       [1:0]    resultStage_controlPipeBeforePipe_s2mPipe_payload_nextPosition;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_horizontalDirectionValid;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_verticalDirectionValid;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_mainDirectionValid;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_counterDirectionValid;
  wire                resultStage_controlPipeBeforePipe_s2mPipe_payload_inValidMinDiff;
  reg                 resultStage_controlPipeBeforePipe_rValid;
  reg                 resultStage_controlPipeBeforePipe_rData_frameStart;
  reg                 resultStage_controlPipeBeforePipe_rData_rowEnd;
  reg                 resultStage_controlPipeBeforePipe_rData_pipeValid;
  reg                 resultStage_controlPipeBeforePipe_rData_firstRow;
  reg                 resultStage_controlPipeBeforePipe_rData_lastRow;
  reg                 resultStage_controlPipeBeforePipe_rData_finalResult;
  reg                 resultStage_controlPipeBeforePipe_rData_mainCompare;
  reg                 resultStage_controlPipeBeforePipe_rData_counterCompare;
  reg                 resultStage_controlPipeBeforePipe_rData_horizontalCompare;
  reg                 resultStage_controlPipeBeforePipe_rData_verticalCompare;
  reg        [7:0]    resultStage_controlPipeBeforePipe_rData_mainDiff;
  reg        [7:0]    resultStage_controlPipeBeforePipe_rData_counterDiff;
  reg        [7:0]    resultStage_controlPipeBeforePipe_rData_horizontalDiff;
  reg        [7:0]    resultStage_controlPipeBeforePipe_rData_verticalDiff;
  reg                 resultStage_controlPipeBeforePipe_rData_isHorizontalMin;
  reg        [7:0]    resultStage_controlPipeBeforePipe_rData_minDiff;
  reg        [1:0]    resultStage_controlPipeBeforePipe_rData_currentPosition;
  reg        [1:0]    resultStage_controlPipeBeforePipe_rData_nextPosition;
  reg                 resultStage_controlPipeBeforePipe_rData_horizontalDirectionValid;
  reg                 resultStage_controlPipeBeforePipe_rData_verticalDirectionValid;
  reg                 resultStage_controlPipeBeforePipe_rData_mainDirectionValid;
  reg                 resultStage_controlPipeBeforePipe_rData_counterDirectionValid;
  reg                 resultStage_controlPipeBeforePipe_rData_inValidMinDiff;
  wire                resultStage_controlPipe_valid;
  wire                resultStage_controlPipe_ready;
  wire                resultStage_controlPipe_payload_frameStart;
  wire                resultStage_controlPipe_payload_rowEnd;
  wire                resultStage_controlPipe_payload_pipeValid;
  wire                resultStage_controlPipe_payload_firstRow;
  wire                resultStage_controlPipe_payload_lastRow;
  wire                resultStage_controlPipe_payload_finalResult;
  wire                resultStage_controlPipe_payload_mainCompare;
  wire                resultStage_controlPipe_payload_counterCompare;
  wire                resultStage_controlPipe_payload_horizontalCompare;
  wire                resultStage_controlPipe_payload_verticalCompare;
  wire       [7:0]    resultStage_controlPipe_payload_mainDiff;
  wire       [7:0]    resultStage_controlPipe_payload_counterDiff;
  wire       [7:0]    resultStage_controlPipe_payload_horizontalDiff;
  wire       [7:0]    resultStage_controlPipe_payload_verticalDiff;
  wire                resultStage_controlPipe_payload_isHorizontalMin;
  wire       [7:0]    resultStage_controlPipe_payload_minDiff;
  wire       [1:0]    resultStage_controlPipe_payload_currentPosition;
  wire       [1:0]    resultStage_controlPipe_payload_nextPosition;
  wire                resultStage_controlPipe_payload_horizontalDirectionValid;
  wire                resultStage_controlPipe_payload_verticalDirectionValid;
  wire                resultStage_controlPipe_payload_mainDirectionValid;
  wire                resultStage_controlPipe_payload_counterDirectionValid;
  wire                resultStage_controlPipe_payload_inValidMinDiff;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rValid;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_frameStart;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_rowEnd;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_pipeValid;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_firstRow;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_lastRow;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_finalResult;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_mainCompare;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_counterCompare;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_horizontalCompare;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_verticalCompare;
  reg        [7:0]    resultStage_controlPipeBeforePipe_s2mPipe_rData_mainDiff;
  reg        [7:0]    resultStage_controlPipeBeforePipe_s2mPipe_rData_counterDiff;
  reg        [7:0]    resultStage_controlPipeBeforePipe_s2mPipe_rData_horizontalDiff;
  reg        [7:0]    resultStage_controlPipeBeforePipe_s2mPipe_rData_verticalDiff;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_isHorizontalMin;
  reg        [7:0]    resultStage_controlPipeBeforePipe_s2mPipe_rData_minDiff;
  reg        [1:0]    resultStage_controlPipeBeforePipe_s2mPipe_rData_currentPosition;
  reg        [1:0]    resultStage_controlPipeBeforePipe_s2mPipe_rData_nextPosition;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_horizontalDirectionValid;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_verticalDirectionValid;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_mainDirectionValid;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_counterDirectionValid;
  reg                 resultStage_controlPipeBeforePipe_s2mPipe_rData_inValidMinDiff;
  wire                when_Stream_l368_66;
  wire                resultStage_pixelStream_valid;
  wire                resultStage_pixelStream_ready;
  reg        [7:0]    resultStage_pixelStream_payload;
  wire                when_SuperResolutionPart3_l840;
  wire                when_SuperResolutionPart3_l846;
  wire                when_SuperResolutionPart3_l847;
  wire                when_SuperResolutionPart3_l850;
  wire                when_SuperResolutionPart3_l854;
  wire                when_SuperResolutionPart3_l855;
  wire                when_SuperResolutionPart3_l860;
  wire                when_SuperResolutionPart3_l861;
  wire                when_SuperResolutionPart3_l851;
  wire                when_SuperResolutionPart3_l841;
  wire                when_SuperResolutionPart3_l842;
  wire                when_SuperResolutionPart3_l869;
  wire                when_SuperResolutionPart3_l870;
  wire                when_SuperResolutionPart3_l871;
  wire                when_SuperResolutionPart3_l872;
  wire                when_SuperResolutionPart3_l875;
  wire                when_SuperResolutionPart3_l876;
  wire                when_SuperResolutionPart3_l885;
  wire                when_SuperResolutionPart3_l893;
  wire                when_SuperResolutionPart3_l884;
  wire                when_SuperResolutionPart3_l902;
  wire                when_SuperResolutionPart3_l903;
  wire                when_SuperResolutionPart3_l912;
  wire                when_SuperResolutionPart3_l920;
  wire                when_SuperResolutionPart3_l911;
  wire                when_SuperResolutionPart3_l874;
  wire                when_SuperResolutionPart3_l930;
  wire                when_SuperResolutionPart3_l931;
  wire                when_SuperResolutionPart3_l932;
  wire                when_SuperResolutionPart3_l941;
  wire                when_SuperResolutionPart3_l949;
  wire                when_SuperResolutionPart3_l940;
  wire                when_SuperResolutionPart3_l958;
  wire                when_SuperResolutionPart3_l959;
  wire                when_SuperResolutionPart3_l968;
  wire                when_SuperResolutionPart3_l976;
  wire                when_SuperResolutionPart3_l967;
  wire                when_SuperResolutionPart3_l986;
  wire                when_SuperResolutionPart3_l987;
  wire                when_SuperResolutionPart3_l988;
  wire                when_SuperResolutionPart3_l991;
  wire                when_SuperResolutionPart3_l992;
  wire                when_SuperResolutionPart3_l1001;
  wire                when_SuperResolutionPart3_l1009;
  wire                when_SuperResolutionPart3_l1000;
  wire                when_SuperResolutionPart3_l1019;
  wire                when_SuperResolutionPart3_l1020;
  wire                when_SuperResolutionPart3_l1021;
  wire                when_SuperResolutionPart3_l1024;
  wire                when_SuperResolutionPart3_l1025;
  wire                when_SuperResolutionPart3_l1034;
  wire                when_SuperResolutionPart3_l1042;
  wire                when_SuperResolutionPart3_l1033;
  wire                when_SuperResolutionPart3_l1052;
  wire                when_SuperResolutionPart3_l1053;
  wire                when_SuperResolutionPart3_l1062;
  wire                when_SuperResolutionPart3_l1070;
  wire                when_SuperResolutionPart3_l1061;
  wire                when_SuperResolutionPart3_l1079;
  wire                when_SuperResolutionPart3_l1080;
  wire                when_SuperResolutionPart3_l1083;
  wire                when_SuperResolutionPart3_l1084;
  wire                when_SuperResolutionPart3_l1093;
  wire                when_SuperResolutionPart3_l1101;
  wire                when_SuperResolutionPart3_l1092;
  wire                when_SuperResolutionPart3_l929;
  wire                when_SuperResolutionPart3_l985;
  wire                when_SuperResolutionPart3_l1018;
  wire                when_SuperResolutionPart3_l1051;
  wire                when_SuperResolutionPart3_l1078;
  wire                when_SuperResolutionPart3_l1082;
  wire                resultStage_pixelStream_s2mPipe_valid;
  reg                 resultStage_pixelStream_s2mPipe_ready;
  wire       [7:0]    resultStage_pixelStream_s2mPipe_payload;
  reg                 resultStage_pixelStream_rValid;
  reg        [7:0]    resultStage_pixelStream_rData;
  wire                resultStage_resultStream_valid;
  wire                resultStage_resultStream_ready;
  wire       [7:0]    resultStage_resultStream_payload;
  reg                 resultStage_pixelStream_s2mPipe_rValid;
  reg        [7:0]    resultStage_pixelStream_s2mPipe_rData;
  wire                when_Stream_l368_67;
  wire                when_SuperResolutionPart3_l1115;
  wire                diffStage_controlPipe_fire;
  wire                CICC1851_resultStage_mainOnePixelStream_ready;
  reg                 CICC1851_resultStage_mainOnePixelStream_ready_1;
  wire                CICC1851_resultStage_mainOnePixelStream_ready_2;
  wire                when_Stream_l438;
  reg                 resultsJoin_valid;
  wire                resultsJoin_ready;
  wire                pixelsStream_valid;
  wire                pixelsStream_ready;
  wire       [7:0]    pixelsStream_payload_pixel;
  wire                pixelsStream_payload_frameStart;
  wire                pixelsStream_payload_rowEnd;
  wire                pixelsStream_s2mPipe_valid;
  reg                 pixelsStream_s2mPipe_ready;
  wire       [7:0]    pixelsStream_s2mPipe_payload_pixel;
  wire                pixelsStream_s2mPipe_payload_frameStart;
  wire                pixelsStream_s2mPipe_payload_rowEnd;
  reg                 pixelsStream_rValid;
  reg        [7:0]    pixelsStream_rData_pixel;
  reg                 pixelsStream_rData_frameStart;
  reg                 pixelsStream_rData_rowEnd;
  wire                pixelsStream_s2mPipe_m2sPipe_valid;
  wire                pixelsStream_s2mPipe_m2sPipe_ready;
  wire       [7:0]    pixelsStream_s2mPipe_m2sPipe_payload_pixel;
  wire                pixelsStream_s2mPipe_m2sPipe_payload_frameStart;
  wire                pixelsStream_s2mPipe_m2sPipe_payload_rowEnd;
  reg                 pixelsStream_s2mPipe_rValid;
  reg        [7:0]    pixelsStream_s2mPipe_rData_pixel;
  reg                 pixelsStream_s2mPipe_rData_frameStart;
  reg                 pixelsStream_s2mPipe_rData_rowEnd;
  wire                when_Stream_l368_68;
  wire                controlStateMachine_wantExit;
  reg                 controlStateMachine_wantStart;
  wire                controlStateMachine_wantKill;
  reg        [1:0]    controlStateMachine_stateReg;
  reg        [1:0]    controlStateMachine_stateNext;
  wire                passPixels_fire_13;
  wire                when_SuperResolutionPart3_l1158;
  wire                controlStream_fire;
  wire                when_SuperResolutionPart3_l1168;
  wire                when_SuperResolutionPart3_l1188;
  wire                controlStream_fire_1;
  wire                when_SuperResolutionPart3_l1199;
  wire                passPixels_fire_14;
  wire                when_SuperResolutionPart3_l1202;
  wire                passPixels_fire_15;
  wire                when_SuperResolutionPart3_l1205;
  wire                when_SuperResolutionPart3_l1217;
  wire                controlStream_fire_2;
  wire                when_SuperResolutionPart3_l1220;
  wire                controlStream_fire_3;
  wire                when_SuperResolutionPart3_l1223;
  wire                controlStream_fire_4;
  wire                when_SuperResolutionPart3_l1224;
  wire                controlStream_fire_5;
  wire                when_SuperResolutionPart3_l1226;
  wire                controlStream_fire_6;
  wire                controlStream_fire_7;
  wire                when_SuperResolutionPart3_l1247;
  wire                when_SuperResolutionPart3_l1248;
  wire                when_SuperResolutionPart3_l1250;
  wire                when_SuperResolutionPart3_l1252;
  `ifndef SYNTHESIS
  reg [39:0] controlStateMachine_stateReg_string;
  reg [39:0] controlStateMachine_stateNext_string;
  `endif

  reg [7:0] lineBufferOne [0:3839];
  reg [7:0] lineBufferTwo [0:3839];
  reg [7:0] lineBufferThree [0:3839];
  reg [0:0] validBufferOne [0:3839];
  reg [0:0] validBufferTwo [0:3839];
  reg [0:0] validBufferThree [0:3839];

  assign CICC1851_bufferRowCount_valueNext_1 = bufferRowCount_willIncrement;
  assign CICC1851_bufferRowCount_valueNext = {11'd0, CICC1851_bufferRowCount_valueNext_1};
  assign CICC1851_bufferWAddr_valueNext_1 = bufferWAddr_willIncrement;
  assign CICC1851_bufferWAddr_valueNext = {11'd0, CICC1851_bufferWAddr_valueNext_1};
  assign CICC1851_outPixelAddr_valueNext_1 = outPixelAddr_willIncrement;
  assign CICC1851_outPixelAddr_valueNext = {11'd0, CICC1851_outPixelAddr_valueNext_1};
  assign CICC1851_outRowCount_valueNext_1 = outRowCount_willIncrement;
  assign CICC1851_outRowCount_valueNext = {11'd0, CICC1851_outRowCount_valueNext_1};
  assign CICC1851_alreadySendRow_valueNext_1 = alreadySendRow_willIncrement;
  assign CICC1851_alreadySendRow_valueNext = {11'd0, CICC1851_alreadySendRow_valueNext_1};
  assign CICC1851_alreadySendCountInRow_valueNext_1 = alreadySendCountInRow_willIncrement;
  assign CICC1851_alreadySendCountInRow_valueNext = {11'd0, CICC1851_alreadySendCountInRow_valueNext_1};
  assign CICC1851_nextRowBuffer = 1'b1;
  assign CICC1851_when_SuperResolutionPart3_l226 = {1'd0, bufferWAddr_value};
  assign CICC1851_when_SuperResolutionPart3_l226_1 = (CICC1851_when_SuperResolutionPart3_l226_2 - 13'h0002);
  assign CICC1851_when_SuperResolutionPart3_l226_2 = (3'b100 * bmpWidth);
  assign CICC1851_when_SuperResolutionPart3_l227 = {1'd0, bufferRowCount_value};
  assign CICC1851_when_SuperResolutionPart3_l227_1 = (CICC1851_when_SuperResolutionPart3_l227_2 - 13'h0002);
  assign CICC1851_when_SuperResolutionPart3_l227_2 = (3'b100 * bmpHeight);
  assign CICC1851_when_SuperResolutionPart3_l270 = {1'd0, alreadySendCountInRow_value};
  assign CICC1851_when_SuperResolutionPart3_l270_1 = (CICC1851_when_SuperResolutionPart3_l270_2 - 13'h0002);
  assign CICC1851_when_SuperResolutionPart3_l270_2 = (3'b100 * bmpWidth);
  assign CICC1851_when_SuperResolutionPart3_l271 = {1'd0, alreadySendRow_value};
  assign CICC1851_when_SuperResolutionPart3_l271_1 = (CICC1851_when_SuperResolutionPart3_l271_2 - 13'h0002);
  assign CICC1851_when_SuperResolutionPart3_l271_2 = (3'b100 * bmpHeight);
  assign CICC1851_resultStage_pixelStream_payload = (CICC1851_resultStage_pixelStream_payload_1 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_1 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_mainThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_2 = (CICC1851_resultStage_pixelStream_payload_3 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_3 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_mainThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_4 = (CICC1851_resultStage_pixelStream_payload_5 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_5 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_mainTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_6 = (CICC1851_resultStage_pixelStream_payload_7 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_7 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_mainThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_8 = (CICC1851_resultStage_pixelStream_payload_9 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_9 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_mainThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_10 = (CICC1851_resultStage_pixelStream_payload_11 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_11 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_mainTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_12 = (CICC1851_resultStage_pixelStream_payload_13 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_13 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_mainThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_14 = (CICC1851_resultStage_pixelStream_payload_15 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_15 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_mainThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_16 = (CICC1851_resultStage_pixelStream_payload_17 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_17 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_mainTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_18 = (CICC1851_resultStage_pixelStream_payload_19 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_19 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_20 = (CICC1851_resultStage_pixelStream_payload_21 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_21 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_22 = (CICC1851_resultStage_pixelStream_payload_23 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_23 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_24 = (CICC1851_resultStage_pixelStream_payload_25 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_25 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_26 = (CICC1851_resultStage_pixelStream_payload_27 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_27 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_28 = (CICC1851_resultStage_pixelStream_payload_29 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_29 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_30 = (CICC1851_resultStage_pixelStream_payload_31 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_31 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_32 = (CICC1851_resultStage_pixelStream_payload_33 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_33 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_34 = (CICC1851_resultStage_pixelStream_payload_35 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_35 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_36 = (CICC1851_resultStage_pixelStream_payload_37 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_37 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_38 = (CICC1851_resultStage_pixelStream_payload_39 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_39 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_40 = (CICC1851_resultStage_pixelStream_payload_41 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_41 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_42 = (CICC1851_resultStage_pixelStream_payload_43 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_43 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_44 = (CICC1851_resultStage_pixelStream_payload_45 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_45 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_46 = (CICC1851_resultStage_pixelStream_payload_47 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_47 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_48 = (CICC1851_resultStage_pixelStream_payload_49 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_49 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_50 = (CICC1851_resultStage_pixelStream_payload_51 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_51 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_52 = (CICC1851_resultStage_pixelStream_payload_53 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_53 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_54 = (CICC1851_resultStage_pixelStream_payload_55 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_55 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_56 = (CICC1851_resultStage_pixelStream_payload_57 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_57 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_58 = (CICC1851_resultStage_pixelStream_payload_59 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_59 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_60 = (CICC1851_resultStage_pixelStream_payload_61 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_61 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_62 = (CICC1851_resultStage_pixelStream_payload_63 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_63 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_64 = (CICC1851_resultStage_pixelStream_payload_65 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_65 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_66 = (CICC1851_resultStage_pixelStream_payload_67 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_67 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_68 = (CICC1851_resultStage_pixelStream_payload_69 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_69 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_70 = (CICC1851_resultStage_pixelStream_payload_71 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_71 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_72 = (CICC1851_resultStage_pixelStream_payload_73 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_73 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_74 = (CICC1851_resultStage_pixelStream_payload_75 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_75 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_76 = (CICC1851_resultStage_pixelStream_payload_77 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_77 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_78 = (CICC1851_resultStage_pixelStream_payload_79 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_79 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_80 = (CICC1851_resultStage_pixelStream_payload_81 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_81 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_82 = (CICC1851_resultStage_pixelStream_payload_83 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_83 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_84 = (CICC1851_resultStage_pixelStream_payload_85 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_85 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_86 = (CICC1851_resultStage_pixelStream_payload_87 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_87 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_88 = (CICC1851_resultStage_pixelStream_payload_89 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_89 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_90 = (CICC1851_resultStage_pixelStream_payload_91 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_91 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_92 = (CICC1851_resultStage_pixelStream_payload_93 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_93 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_94 = (CICC1851_resultStage_pixelStream_payload_95 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_95 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_96 = (CICC1851_resultStage_pixelStream_payload_97 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_97 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_98 = (CICC1851_resultStage_pixelStream_payload_99 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_99 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_100 = (CICC1851_resultStage_pixelStream_payload_101 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_101 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_102 = (CICC1851_resultStage_pixelStream_payload_103 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_103 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_104 = (CICC1851_resultStage_pixelStream_payload_105 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_105 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_106 = (CICC1851_resultStage_pixelStream_payload_107 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_107 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_108 = (CICC1851_resultStage_pixelStream_payload_109 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_109 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_110 = (CICC1851_resultStage_pixelStream_payload_111 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_111 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_112 = (CICC1851_resultStage_pixelStream_payload_113 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_113 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_114 = (CICC1851_resultStage_pixelStream_payload_115 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_115 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_116 = (CICC1851_resultStage_pixelStream_payload_117 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_117 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_118 = (CICC1851_resultStage_pixelStream_payload_119 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_119 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_120 = (CICC1851_resultStage_pixelStream_payload_121 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_121 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_122 = (CICC1851_resultStage_pixelStream_payload_123 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_123 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_124 = (CICC1851_resultStage_pixelStream_payload_125 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_125 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_126 = (CICC1851_resultStage_pixelStream_payload_127 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_127 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_128 = (CICC1851_resultStage_pixelStream_payload_129 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_129 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_130 = (CICC1851_resultStage_pixelStream_payload_131 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_131 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_132 = (CICC1851_resultStage_pixelStream_payload_133 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_133 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_134 = (CICC1851_resultStage_pixelStream_payload_135 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_135 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_136 = (CICC1851_resultStage_pixelStream_payload_137 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_137 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_138 = (CICC1851_resultStage_pixelStream_payload_139 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_139 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_140 = (CICC1851_resultStage_pixelStream_payload_141 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_141 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_142 = (CICC1851_resultStage_pixelStream_payload_143 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_143 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_144 = (CICC1851_resultStage_pixelStream_payload_145 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_145 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_146 = (CICC1851_resultStage_pixelStream_payload_147 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_147 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_148 = (CICC1851_resultStage_pixelStream_payload_149 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_149 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_150 = (CICC1851_resultStage_pixelStream_payload_151 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_151 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_152 = (CICC1851_resultStage_pixelStream_payload_153 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_153 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_154 = (CICC1851_resultStage_pixelStream_payload_155 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_155 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_156 = (CICC1851_resultStage_pixelStream_payload_157 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_157 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_158 = (CICC1851_resultStage_pixelStream_payload_159 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_159 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_160 = (CICC1851_resultStage_pixelStream_payload_161 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_161 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_162 = (CICC1851_resultStage_pixelStream_payload_163 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_163 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_164 = (CICC1851_resultStage_pixelStream_payload_165 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_165 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_166 = (CICC1851_resultStage_pixelStream_payload_167 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_167 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_168 = (CICC1851_resultStage_pixelStream_payload_169 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_169 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_170 = (CICC1851_resultStage_pixelStream_payload_171 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_171 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_172 = (CICC1851_resultStage_pixelStream_payload_173 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_173 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_174 = (CICC1851_resultStage_pixelStream_payload_175 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_175 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_176 = (CICC1851_resultStage_pixelStream_payload_177 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_177 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_178 = (CICC1851_resultStage_pixelStream_payload_179 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_179 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_180 = (CICC1851_resultStage_pixelStream_payload_181 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_181 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_182 = (CICC1851_resultStage_pixelStream_payload_183 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_183 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_184 = (CICC1851_resultStage_pixelStream_payload_185 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_185 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_186 = (CICC1851_resultStage_pixelStream_payload_187 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_187 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_188 = (CICC1851_resultStage_pixelStream_payload_189 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_189 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_190 = (CICC1851_resultStage_pixelStream_payload_191 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_191 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_192 = (CICC1851_resultStage_pixelStream_payload_193 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_193 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_194 = (CICC1851_resultStage_pixelStream_payload_195 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_195 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_196 = (CICC1851_resultStage_pixelStream_payload_197 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_197 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_198 = (CICC1851_resultStage_pixelStream_payload_199 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_199 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_200 = (CICC1851_resultStage_pixelStream_payload_201 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_201 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_202 = (CICC1851_resultStage_pixelStream_payload_203 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_203 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_204 = (CICC1851_resultStage_pixelStream_payload_205 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_205 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_206 = (CICC1851_resultStage_pixelStream_payload_207 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_207 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_208 = (CICC1851_resultStage_pixelStream_payload_209 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_209 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_210 = (CICC1851_resultStage_pixelStream_payload_211 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_211 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_212 = (CICC1851_resultStage_pixelStream_payload_213 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_213 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_214 = (CICC1851_resultStage_pixelStream_payload_215 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_215 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_216 = (CICC1851_resultStage_pixelStream_payload_217 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_217 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_218 = (CICC1851_resultStage_pixelStream_payload_219 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_219 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_220 = (CICC1851_resultStage_pixelStream_payload_221 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_221 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_222 = (CICC1851_resultStage_pixelStream_payload_223 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_223 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_224 = (CICC1851_resultStage_pixelStream_payload_225 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_225 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_226 = (CICC1851_resultStage_pixelStream_payload_227 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_227 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_228 = (CICC1851_resultStage_pixelStream_payload_229 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_229 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_230 = (CICC1851_resultStage_pixelStream_payload_231 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_231 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_232 = (CICC1851_resultStage_pixelStream_payload_233 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_233 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_234 = (CICC1851_resultStage_pixelStream_payload_235 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_235 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_236 = (CICC1851_resultStage_pixelStream_payload_237 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_237 = ({1'b0,diffStage_mainThreePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_238 = (CICC1851_resultStage_pixelStream_payload_239 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_239 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_240 = (CICC1851_resultStage_pixelStream_payload_241 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_241 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterThreePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_242 = (CICC1851_resultStage_pixelStream_payload_243 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_243 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_244 = (CICC1851_resultStage_pixelStream_payload_245 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_245 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_246 = (CICC1851_resultStage_pixelStream_payload_247 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_247 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_248 = (CICC1851_resultStage_pixelStream_payload_249 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_249 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_when_SuperResolutionPart3_l1202 = (12'h003 + outRowCount_value);
  assign CICC1851_when_SuperResolutionPart3_l1205 = (12'h001 + outRowCount_value);
  assign CICC1851_when_SuperResolutionPart3_l1205_1 = (12'h002 + outPixelAddr_value);
  assign CICC1851_when_SuperResolutionPart3_l1205_2 = (12'h002 + outPixelAddr_value);
  assign CICC1851_when_SuperResolutionPart3_l1223 = {1'd0, outPixelAddr_value};
  assign CICC1851_when_SuperResolutionPart3_l1223_1 = (CICC1851_when_SuperResolutionPart3_l1223_2 - 13'h0002);
  assign CICC1851_when_SuperResolutionPart3_l1223_2 = (3'b100 * bmpWidth);
  assign CICC1851_when_SuperResolutionPart3_l1224 = {1'd0, outRowCount_value};
  assign CICC1851_when_SuperResolutionPart3_l1224_1 = (CICC1851_when_SuperResolutionPart3_l1224_2 - 13'h0002);
  assign CICC1851_when_SuperResolutionPart3_l1224_2 = (3'b100 * bmpHeight);
  assign CICC1851_lineBufferOne_port = passPixels_payload_pixel;
  assign CICC1851_lineBufferOne_port_1 = (passPixels_fire_6 && (bufferSwitch == 2'b00));
  assign CICC1851_lineBufferTwo_port = passPixels_payload_pixel;
  assign CICC1851_lineBufferTwo_port_1 = (passPixels_fire_7 && (bufferSwitch == 2'b01));
  assign CICC1851_lineBufferThree_port = passPixels_payload_pixel;
  assign CICC1851_lineBufferThree_port_1 = (passPixels_fire_8 && (bufferSwitch == 2'b10));
  assign CICC1851_validBufferOne_port = passPixels_payload_inpValid;
  assign CICC1851_validBufferOne_port_1 = (passPixels_fire_9 && (bufferSwitch == 2'b00));
  assign CICC1851_validBufferTwo_port = passPixels_payload_inpValid;
  assign CICC1851_validBufferTwo_port_1 = (passPixels_fire_10 && (bufferSwitch == 2'b01));
  assign CICC1851_validBufferThree_port = passPixels_payload_inpValid;
  assign CICC1851_validBufferThree_port_1 = (passPixels_fire_11 && (bufferSwitch == 2'b10));
  always @(posedge clk) begin
    if(CICC1851_lineBufferOne_port_1) begin
      lineBufferOne[bufferWAddr_value] <= CICC1851_lineBufferOne_port;
    end
  end

  always @(posedge clk) begin
    if(mainPixelAddrOneStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferOne_port1 <= lineBufferOne[mainPixelAddrOneStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(counterPixelAddrOneStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferOne_port2 <= lineBufferOne[counterPixelAddrOneStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(CICC1851_lineBufferTwo_port_1) begin
      lineBufferTwo[bufferWAddr_value] <= CICC1851_lineBufferTwo_port;
    end
  end

  always @(posedge clk) begin
    if(mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferTwo_port1 <= lineBufferTwo[mainPixelAddrTwoStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferTwo_port2 <= lineBufferTwo[counterPixelAddrTwoStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(CICC1851_lineBufferThree_port_1) begin
      lineBufferThree[bufferWAddr_value] <= CICC1851_lineBufferThree_port;
    end
  end

  always @(posedge clk) begin
    if(mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferThree_port1 <= lineBufferThree[mainPixelAddrThreeStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferThree_port2 <= lineBufferThree[counterPixelAddrThreeStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(CICC1851_validBufferOne_port_1) begin
      validBufferOne[bufferWAddr_value] <= CICC1851_validBufferOne_port;
    end
  end

  always @(posedge clk) begin
    if(mainValidAddrOneStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_validBufferOne_port1 <= validBufferOne[mainValidAddrOneStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(counterValidAddrOneStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_validBufferOne_port2 <= validBufferOne[counterValidAddrOneStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(CICC1851_validBufferTwo_port_1) begin
      validBufferTwo[bufferWAddr_value] <= CICC1851_validBufferTwo_port;
    end
  end

  always @(posedge clk) begin
    if(mainValidAddrTwoStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_validBufferTwo_port1 <= validBufferTwo[mainValidAddrTwoStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(counterValidAddrTwoStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_validBufferTwo_port2 <= validBufferTwo[counterValidAddrTwoStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(CICC1851_validBufferThree_port_1) begin
      validBufferThree[bufferWAddr_value] <= CICC1851_validBufferThree_port;
    end
  end

  always @(posedge clk) begin
    if(mainValidAddrThreeStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_validBufferThree_port1 <= validBufferThree[mainValidAddrThreeStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(counterValidAddrThreeStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_validBufferThree_port2 <= validBufferThree[counterValidAddrThreeStream_s2mPipe_m2sPipe_payload];
    end
  end

  StreamFork_3 diffStage_controlPipe_fork (
    .io_input_valid                                (diffStage_controlPipe_valid                                             ), //i
    .io_input_ready                                (diffStage_controlPipe_fork_io_input_ready                               ), //o
    .io_input_payload_frameStart                   (diffStage_controlPipe_payload_frameStart                                ), //i
    .io_input_payload_rowEnd                       (diffStage_controlPipe_payload_rowEnd                                    ), //i
    .io_input_payload_pipeValid                    (diffStage_controlPipe_payload_pipeValid                                 ), //i
    .io_input_payload_firstRow                     (diffStage_controlPipe_payload_firstRow                                  ), //i
    .io_input_payload_lastRow                      (diffStage_controlPipe_payload_lastRow                                   ), //i
    .io_input_payload_finalResult                  (diffStage_controlPipe_payload_finalResult                               ), //i
    .io_input_payload_mainCompare                  (diffStage_controlPipe_payload_mainCompare                               ), //i
    .io_input_payload_counterCompare               (diffStage_controlPipe_payload_counterCompare                            ), //i
    .io_input_payload_horizontalCompare            (diffStage_controlPipe_payload_horizontalCompare                         ), //i
    .io_input_payload_verticalCompare              (diffStage_controlPipe_payload_verticalCompare                           ), //i
    .io_input_payload_mainDiff                     (diffStage_controlPipe_payload_mainDiff[7:0]                             ), //i
    .io_input_payload_counterDiff                  (diffStage_controlPipe_payload_counterDiff[7:0]                          ), //i
    .io_input_payload_horizontalDiff               (diffStage_controlPipe_payload_horizontalDiff[7:0]                       ), //i
    .io_input_payload_verticalDiff                 (diffStage_controlPipe_payload_verticalDiff[7:0]                         ), //i
    .io_input_payload_isHorizontalMin              (diffStage_controlPipe_payload_isHorizontalMin                           ), //i
    .io_input_payload_minDiff                      (diffStage_controlPipe_payload_minDiff[7:0]                              ), //i
    .io_input_payload_currentPosition              (diffStage_controlPipe_payload_currentPosition[1:0]                      ), //i
    .io_input_payload_nextPosition                 (diffStage_controlPipe_payload_nextPosition[1:0]                         ), //i
    .io_input_payload_horizontalDirectionValid     (diffStage_controlPipe_payload_horizontalDirectionValid                  ), //i
    .io_input_payload_verticalDirectionValid       (diffStage_controlPipe_payload_verticalDirectionValid                    ), //i
    .io_input_payload_mainDirectionValid           (diffStage_controlPipe_payload_mainDirectionValid                        ), //i
    .io_input_payload_counterDirectionValid        (diffStage_controlPipe_payload_counterDirectionValid                     ), //i
    .io_input_payload_inValidMinDiff               (diffStage_controlPipe_payload_inValidMinDiff                            ), //i
    .io_outputs_0_valid                            (diffStage_controlPipe_fork_io_outputs_0_valid                           ), //o
    .io_outputs_0_ready                            (resultStage_controlPipeBeforePipe_ready                                 ), //i
    .io_outputs_0_payload_frameStart               (diffStage_controlPipe_fork_io_outputs_0_payload_frameStart              ), //o
    .io_outputs_0_payload_rowEnd                   (diffStage_controlPipe_fork_io_outputs_0_payload_rowEnd                  ), //o
    .io_outputs_0_payload_pipeValid                (diffStage_controlPipe_fork_io_outputs_0_payload_pipeValid               ), //o
    .io_outputs_0_payload_firstRow                 (diffStage_controlPipe_fork_io_outputs_0_payload_firstRow                ), //o
    .io_outputs_0_payload_lastRow                  (diffStage_controlPipe_fork_io_outputs_0_payload_lastRow                 ), //o
    .io_outputs_0_payload_finalResult              (diffStage_controlPipe_fork_io_outputs_0_payload_finalResult             ), //o
    .io_outputs_0_payload_mainCompare              (diffStage_controlPipe_fork_io_outputs_0_payload_mainCompare             ), //o
    .io_outputs_0_payload_counterCompare           (diffStage_controlPipe_fork_io_outputs_0_payload_counterCompare          ), //o
    .io_outputs_0_payload_horizontalCompare        (diffStage_controlPipe_fork_io_outputs_0_payload_horizontalCompare       ), //o
    .io_outputs_0_payload_verticalCompare          (diffStage_controlPipe_fork_io_outputs_0_payload_verticalCompare         ), //o
    .io_outputs_0_payload_mainDiff                 (diffStage_controlPipe_fork_io_outputs_0_payload_mainDiff[7:0]           ), //o
    .io_outputs_0_payload_counterDiff              (diffStage_controlPipe_fork_io_outputs_0_payload_counterDiff[7:0]        ), //o
    .io_outputs_0_payload_horizontalDiff           (diffStage_controlPipe_fork_io_outputs_0_payload_horizontalDiff[7:0]     ), //o
    .io_outputs_0_payload_verticalDiff             (diffStage_controlPipe_fork_io_outputs_0_payload_verticalDiff[7:0]       ), //o
    .io_outputs_0_payload_isHorizontalMin          (diffStage_controlPipe_fork_io_outputs_0_payload_isHorizontalMin         ), //o
    .io_outputs_0_payload_minDiff                  (diffStage_controlPipe_fork_io_outputs_0_payload_minDiff[7:0]            ), //o
    .io_outputs_0_payload_currentPosition          (diffStage_controlPipe_fork_io_outputs_0_payload_currentPosition[1:0]    ), //o
    .io_outputs_0_payload_nextPosition             (diffStage_controlPipe_fork_io_outputs_0_payload_nextPosition[1:0]       ), //o
    .io_outputs_0_payload_horizontalDirectionValid (diffStage_controlPipe_fork_io_outputs_0_payload_horizontalDirectionValid), //o
    .io_outputs_0_payload_verticalDirectionValid   (diffStage_controlPipe_fork_io_outputs_0_payload_verticalDirectionValid  ), //o
    .io_outputs_0_payload_mainDirectionValid       (diffStage_controlPipe_fork_io_outputs_0_payload_mainDirectionValid      ), //o
    .io_outputs_0_payload_counterDirectionValid    (diffStage_controlPipe_fork_io_outputs_0_payload_counterDirectionValid   ), //o
    .io_outputs_0_payload_inValidMinDiff           (diffStage_controlPipe_fork_io_outputs_0_payload_inValidMinDiff          ), //o
    .io_outputs_1_valid                            (diffStage_controlPipe_fork_io_outputs_1_valid                           ), //o
    .io_outputs_1_ready                            (resultStage_pixelStream_ready                                           ), //i
    .io_outputs_1_payload_frameStart               (diffStage_controlPipe_fork_io_outputs_1_payload_frameStart              ), //o
    .io_outputs_1_payload_rowEnd                   (diffStage_controlPipe_fork_io_outputs_1_payload_rowEnd                  ), //o
    .io_outputs_1_payload_pipeValid                (diffStage_controlPipe_fork_io_outputs_1_payload_pipeValid               ), //o
    .io_outputs_1_payload_firstRow                 (diffStage_controlPipe_fork_io_outputs_1_payload_firstRow                ), //o
    .io_outputs_1_payload_lastRow                  (diffStage_controlPipe_fork_io_outputs_1_payload_lastRow                 ), //o
    .io_outputs_1_payload_finalResult              (diffStage_controlPipe_fork_io_outputs_1_payload_finalResult             ), //o
    .io_outputs_1_payload_mainCompare              (diffStage_controlPipe_fork_io_outputs_1_payload_mainCompare             ), //o
    .io_outputs_1_payload_counterCompare           (diffStage_controlPipe_fork_io_outputs_1_payload_counterCompare          ), //o
    .io_outputs_1_payload_horizontalCompare        (diffStage_controlPipe_fork_io_outputs_1_payload_horizontalCompare       ), //o
    .io_outputs_1_payload_verticalCompare          (diffStage_controlPipe_fork_io_outputs_1_payload_verticalCompare         ), //o
    .io_outputs_1_payload_mainDiff                 (diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff[7:0]           ), //o
    .io_outputs_1_payload_counterDiff              (diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff[7:0]        ), //o
    .io_outputs_1_payload_horizontalDiff           (diffStage_controlPipe_fork_io_outputs_1_payload_horizontalDiff[7:0]     ), //o
    .io_outputs_1_payload_verticalDiff             (diffStage_controlPipe_fork_io_outputs_1_payload_verticalDiff[7:0]       ), //o
    .io_outputs_1_payload_isHorizontalMin          (diffStage_controlPipe_fork_io_outputs_1_payload_isHorizontalMin         ), //o
    .io_outputs_1_payload_minDiff                  (diffStage_controlPipe_fork_io_outputs_1_payload_minDiff[7:0]            ), //o
    .io_outputs_1_payload_currentPosition          (diffStage_controlPipe_fork_io_outputs_1_payload_currentPosition[1:0]    ), //o
    .io_outputs_1_payload_nextPosition             (diffStage_controlPipe_fork_io_outputs_1_payload_nextPosition[1:0]       ), //o
    .io_outputs_1_payload_horizontalDirectionValid (diffStage_controlPipe_fork_io_outputs_1_payload_horizontalDirectionValid), //o
    .io_outputs_1_payload_verticalDirectionValid   (diffStage_controlPipe_fork_io_outputs_1_payload_verticalDirectionValid  ), //o
    .io_outputs_1_payload_mainDirectionValid       (diffStage_controlPipe_fork_io_outputs_1_payload_mainDirectionValid      ), //o
    .io_outputs_1_payload_counterDirectionValid    (diffStage_controlPipe_fork_io_outputs_1_payload_counterDirectionValid   ), //o
    .io_outputs_1_payload_inValidMinDiff           (diffStage_controlPipe_fork_io_outputs_1_payload_inValidMinDiff          )  //o
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_2_BOOT : controlStateMachine_stateReg_string = "BOOT ";
      controlStateMachine_enumDef_2_HOLD : controlStateMachine_stateReg_string = "HOLD ";
      controlStateMachine_enumDef_2_PASS : controlStateMachine_stateReg_string = "PASS ";
      controlStateMachine_enumDef_2_EXTRA : controlStateMachine_stateReg_string = "EXTRA";
      default : controlStateMachine_stateReg_string = "?????";
    endcase
  end
  always @(*) begin
    case(controlStateMachine_stateNext)
      controlStateMachine_enumDef_2_BOOT : controlStateMachine_stateNext_string = "BOOT ";
      controlStateMachine_enumDef_2_HOLD : controlStateMachine_stateNext_string = "HOLD ";
      controlStateMachine_enumDef_2_PASS : controlStateMachine_stateNext_string = "PASS ";
      controlStateMachine_enumDef_2_EXTRA : controlStateMachine_stateNext_string = "EXTRA";
      default : controlStateMachine_stateNext_string = "?????";
    endcase
  end
  `endif

  always @(*) begin
    pixelsIn_ready = 1'b0;
    pixelsIn_ready = (! pixelsIn_rValid);
  end

  always @(*) begin
    pixelsOut_valid = 1'b0;
    pixelsOut_valid = pixelsStream_s2mPipe_m2sPipe_valid;
  end

  always @(*) begin
    pixelsOut_payload_pixel = 8'h0;
    pixelsOut_payload_pixel = pixelsStream_s2mPipe_m2sPipe_payload_pixel;
  end

  always @(*) begin
    pixelsOut_payload_frameStart = 1'b0;
    pixelsOut_payload_frameStart = pixelsStream_s2mPipe_m2sPipe_payload_frameStart;
  end

  always @(*) begin
    pixelsOut_payload_rowEnd = 1'b0;
    pixelsOut_payload_rowEnd = pixelsStream_s2mPipe_m2sPipe_payload_rowEnd;
  end

  always @(*) begin
    inpThreeDoneOut = 1'b0;
    inpThreeDoneOut = inpThreeDone;
  end

  assign when_SuperResolutionPart3_l72 = (startIn && (! startIn_regNext));
  assign when_SuperResolutionPart3_l75 = (! startIn);
  assign when_SuperResolutionPart3_l78 = (startIn && (! readDone));
  assign when_SuperResolutionPart3_l78_1 = (! startIn);
  assign when_SuperResolutionPart3_l93 = (! startIn);
  assign when_SuperResolutionPart3_l96 = (! startIn);
  always @(*) begin
    bufferRowCount_willIncrement = 1'b0;
    if(when_SuperResolutionPart3_l230) begin
      if(!bufferReachFinalRow) begin
        bufferRowCount_willIncrement = 1'b1;
      end
    end
  end

  always @(*) begin
    bufferRowCount_willClear = 1'b0;
    if(when_SuperResolutionPart3_l230) begin
      if(bufferReachFinalRow) begin
        bufferRowCount_willClear = 1'b1;
      end
    end
  end

  assign bufferRowCount_willOverflowIfInc = (bufferRowCount_value == 12'h870);
  assign bufferRowCount_willOverflow = (bufferRowCount_willOverflowIfInc && bufferRowCount_willIncrement);
  always @(*) begin
    if(bufferRowCount_willOverflow) begin
      bufferRowCount_valueNext = 12'h0;
    end else begin
      bufferRowCount_valueNext = (bufferRowCount_value + CICC1851_bufferRowCount_valueNext);
    end
    if(bufferRowCount_willClear) begin
      bufferRowCount_valueNext = 12'h0;
    end
  end

  assign when_SuperResolutionPart3_l102 = ((startIn && (! holdBuffer)) && (! writeDone));
  assign when_SuperResolutionPart3_l102_1 = (((! startIn) || holdBuffer) || writeDone);
  always @(*) begin
    bufferWAddr_willIncrement = 1'b0;
    if(passPixels_fire_12) begin
      if(!passPixels_payload_rowEnd) begin
        bufferWAddr_willIncrement = 1'b1;
      end
    end
  end

  always @(*) begin
    bufferWAddr_willClear = 1'b0;
    if(passPixels_fire_12) begin
      if(passPixels_payload_rowEnd) begin
        bufferWAddr_willClear = 1'b1;
      end
    end
  end

  assign bufferWAddr_willOverflowIfInc = (bufferWAddr_value == 12'heff);
  assign bufferWAddr_willOverflow = (bufferWAddr_willOverflowIfInc && bufferWAddr_willIncrement);
  always @(*) begin
    if(bufferWAddr_willOverflow) begin
      bufferWAddr_valueNext = 12'h0;
    end else begin
      bufferWAddr_valueNext = (bufferWAddr_value + CICC1851_bufferWAddr_valueNext);
    end
    if(bufferWAddr_willClear) begin
      bufferWAddr_valueNext = 12'h0;
    end
  end

  always @(*) begin
    outPixelAddr_willIncrement = 1'b0;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_2_HOLD : begin
      end
      controlStateMachine_enumDef_2_PASS : begin
      end
      controlStateMachine_enumDef_2_EXTRA : begin
        if(controlStream_fire_6) begin
          if(!outReachRowEnd) begin
            outPixelAddr_willIncrement = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outPixelAddr_willClear = 1'b0;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_2_HOLD : begin
      end
      controlStateMachine_enumDef_2_PASS : begin
      end
      controlStateMachine_enumDef_2_EXTRA : begin
        if(controlStream_fire_6) begin
          if(outReachRowEnd) begin
            outPixelAddr_willClear = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign outPixelAddr_willOverflowIfInc = (outPixelAddr_value == 12'heff);
  assign outPixelAddr_willOverflow = (outPixelAddr_willOverflowIfInc && outPixelAddr_willIncrement);
  always @(*) begin
    if(outPixelAddr_willOverflow) begin
      outPixelAddr_valueNext = 12'h0;
    end else begin
      outPixelAddr_valueNext = (outPixelAddr_value + CICC1851_outPixelAddr_valueNext);
    end
    if(outPixelAddr_willClear) begin
      outPixelAddr_valueNext = 12'h0;
    end
  end

  always @(*) begin
    outRowCount_willIncrement = 1'b0;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_2_HOLD : begin
      end
      controlStateMachine_enumDef_2_PASS : begin
      end
      controlStateMachine_enumDef_2_EXTRA : begin
        if(when_SuperResolutionPart3_l1226) begin
          if(!outReachFinalRow) begin
            outRowCount_willIncrement = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outRowCount_willClear = 1'b0;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_2_HOLD : begin
      end
      controlStateMachine_enumDef_2_PASS : begin
      end
      controlStateMachine_enumDef_2_EXTRA : begin
        if(when_SuperResolutionPart3_l1226) begin
          if(outReachFinalRow) begin
            outRowCount_willClear = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign outRowCount_willOverflowIfInc = (outRowCount_value == 12'h870);
  assign outRowCount_willOverflow = (outRowCount_willOverflowIfInc && outRowCount_willIncrement);
  always @(*) begin
    if(outRowCount_willOverflow) begin
      outRowCount_valueNext = 12'h0;
    end else begin
      outRowCount_valueNext = (outRowCount_value + CICC1851_outRowCount_valueNext);
    end
    if(outRowCount_willClear) begin
      outRowCount_valueNext = 12'h0;
    end
  end

  always @(*) begin
    alreadySendRow_willIncrement = 1'b0;
    if(pixelsOut_fire_2) begin
      if(alreadyReachRowEnd) begin
        if(!alreadyReachFinalRow) begin
          alreadySendRow_willIncrement = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    alreadySendRow_willClear = 1'b0;
    if(pixelsOut_fire_2) begin
      if(alreadyReachRowEnd) begin
        if(alreadyReachFinalRow) begin
          alreadySendRow_willClear = 1'b1;
        end
      end
    end
  end

  assign alreadySendRow_willOverflowIfInc = (alreadySendRow_value == 12'h870);
  assign alreadySendRow_willOverflow = (alreadySendRow_willOverflowIfInc && alreadySendRow_willIncrement);
  always @(*) begin
    if(alreadySendRow_willOverflow) begin
      alreadySendRow_valueNext = 12'h0;
    end else begin
      alreadySendRow_valueNext = (alreadySendRow_value + CICC1851_alreadySendRow_valueNext);
    end
    if(alreadySendRow_willClear) begin
      alreadySendRow_valueNext = 12'h0;
    end
  end

  always @(*) begin
    alreadySendCountInRow_willIncrement = 1'b0;
    if(pixelsOut_fire_2) begin
      if(!alreadyReachRowEnd) begin
        alreadySendCountInRow_willIncrement = 1'b1;
      end
    end
  end

  always @(*) begin
    alreadySendCountInRow_willClear = 1'b0;
    if(pixelsOut_fire_2) begin
      if(alreadyReachRowEnd) begin
        alreadySendCountInRow_willClear = 1'b1;
      end
    end
  end

  assign alreadySendCountInRow_willOverflowIfInc = (alreadySendCountInRow_value == 12'heff);
  assign alreadySendCountInRow_willOverflow = (alreadySendCountInRow_willOverflowIfInc && alreadySendCountInRow_willIncrement);
  always @(*) begin
    if(alreadySendCountInRow_willOverflow) begin
      alreadySendCountInRow_valueNext = 12'h0;
    end else begin
      alreadySendCountInRow_valueNext = (alreadySendCountInRow_value + CICC1851_alreadySendCountInRow_valueNext);
    end
    if(alreadySendCountInRow_willClear) begin
      alreadySendCountInRow_valueNext = 12'h0;
    end
  end

  assign when_SuperResolutionPart3_l154 = ((! startRead) || ((! startIn) && startIn_regNext_1));
  always @(*) begin
    mainAddrOne = outPixelAddr_value;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_2_HOLD : begin
      end
      controlStateMachine_enumDef_2_PASS : begin
        if(when_SuperResolutionPart3_l1168) begin
          mainAddrOne = (12'h001 + outPixelAddr_value);
        end else begin
          mainAddrOne = (outPixelAddr_value - 12'h001);
        end
      end
      controlStateMachine_enumDef_2_EXTRA : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    counterAddrOne = outPixelAddr_value;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_2_HOLD : begin
      end
      controlStateMachine_enumDef_2_PASS : begin
        if(outReachRowEnd) begin
          counterAddrOne = (outPixelAddr_value - 12'h001);
        end else begin
          counterAddrOne = (12'h001 + outPixelAddr_value);
        end
      end
      controlStateMachine_enumDef_2_EXTRA : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    mainAddrTwo = outPixelAddr_value;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_2_HOLD : begin
      end
      controlStateMachine_enumDef_2_PASS : begin
        if(when_SuperResolutionPart3_l1168) begin
          mainAddrTwo = (12'h001 + outPixelAddr_value);
        end else begin
          mainAddrTwo = (outPixelAddr_value - 12'h001);
        end
      end
      controlStateMachine_enumDef_2_EXTRA : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    counterAddrTwo = outPixelAddr_value;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_2_HOLD : begin
      end
      controlStateMachine_enumDef_2_PASS : begin
        if(outReachRowEnd) begin
          counterAddrTwo = (outPixelAddr_value - 12'h001);
        end else begin
          counterAddrTwo = (12'h001 + outPixelAddr_value);
        end
      end
      controlStateMachine_enumDef_2_EXTRA : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    mainAddrThree = outPixelAddr_value;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_2_HOLD : begin
      end
      controlStateMachine_enumDef_2_PASS : begin
        if(when_SuperResolutionPart3_l1168) begin
          mainAddrThree = (12'h001 + outPixelAddr_value);
        end else begin
          mainAddrThree = (outPixelAddr_value - 12'h001);
        end
      end
      controlStateMachine_enumDef_2_EXTRA : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    counterAddrThree = outPixelAddr_value;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_2_HOLD : begin
      end
      controlStateMachine_enumDef_2_PASS : begin
        if(outReachRowEnd) begin
          counterAddrThree = (outPixelAddr_value - 12'h001);
        end else begin
          counterAddrThree = (12'h001 + outPixelAddr_value);
        end
      end
      controlStateMachine_enumDef_2_EXTRA : begin
      end
      default : begin
      end
    endcase
  end

  assign validStream_valid = 1'b1;
  assign CICC1851_controls_frameStart = 60'h0;
  always @(*) begin
    controls_frameStart = CICC1851_controls_frameStart[0];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_2_HOLD : begin
      end
      controlStateMachine_enumDef_2_PASS : begin
        if(frameStart) begin
          controls_frameStart = 1'b1;
        end
      end
      controlStateMachine_enumDef_2_EXTRA : begin
        if(frameStart) begin
          controls_frameStart = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_rowEnd = CICC1851_controls_frameStart[1];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_2_HOLD : begin
      end
      controlStateMachine_enumDef_2_PASS : begin
        if(outReachRowEnd) begin
          controls_rowEnd = 1'b1;
        end
      end
      controlStateMachine_enumDef_2_EXTRA : begin
        if(outReachRowEnd) begin
          controls_rowEnd = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_pipeValid = CICC1851_controls_frameStart[2];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_2_HOLD : begin
      end
      controlStateMachine_enumDef_2_PASS : begin
        controls_pipeValid = 1'b1;
      end
      controlStateMachine_enumDef_2_EXTRA : begin
        controls_pipeValid = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_firstRow = CICC1851_controls_frameStart[3];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_2_HOLD : begin
      end
      controlStateMachine_enumDef_2_PASS : begin
        if(when_SuperResolutionPart3_l1188) begin
          controls_firstRow = 1'b1;
        end
      end
      controlStateMachine_enumDef_2_EXTRA : begin
        if(when_SuperResolutionPart3_l1217) begin
          controls_firstRow = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_lastRow = CICC1851_controls_frameStart[4];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_2_HOLD : begin
      end
      controlStateMachine_enumDef_2_PASS : begin
        if(outReachFinalRow) begin
          controls_lastRow = 1'b1;
        end
      end
      controlStateMachine_enumDef_2_EXTRA : begin
        if(outReachFinalRow) begin
          controls_lastRow = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_finalResult = CICC1851_controls_frameStart[5];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_2_HOLD : begin
      end
      controlStateMachine_enumDef_2_PASS : begin
      end
      controlStateMachine_enumDef_2_EXTRA : begin
        controls_finalResult = 1'b1;
      end
      default : begin
      end
    endcase
  end

  assign controls_mainCompare = CICC1851_controls_frameStart[6];
  assign controls_counterCompare = CICC1851_controls_frameStart[7];
  assign controls_horizontalCompare = CICC1851_controls_frameStart[8];
  assign controls_verticalCompare = CICC1851_controls_frameStart[9];
  assign controls_mainDiff = CICC1851_controls_frameStart[17 : 10];
  assign controls_counterDiff = CICC1851_controls_frameStart[25 : 18];
  assign controls_horizontalDiff = CICC1851_controls_frameStart[33 : 26];
  assign controls_verticalDiff = CICC1851_controls_frameStart[41 : 34];
  assign controls_isHorizontalMin = CICC1851_controls_frameStart[42];
  assign controls_minDiff = CICC1851_controls_frameStart[50 : 43];
  always @(*) begin
    controls_currentPosition = CICC1851_controls_frameStart[52 : 51];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_2_HOLD : begin
      end
      controlStateMachine_enumDef_2_PASS : begin
        controls_currentPosition = currentRowBuffer;
      end
      controlStateMachine_enumDef_2_EXTRA : begin
        controls_currentPosition = currentRowBuffer;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_nextPosition = CICC1851_controls_frameStart[54 : 53];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_2_HOLD : begin
      end
      controlStateMachine_enumDef_2_PASS : begin
        controls_nextPosition = nextRowBuffer;
      end
      controlStateMachine_enumDef_2_EXTRA : begin
        controls_nextPosition = nextRowBuffer;
      end
      default : begin
      end
    endcase
  end

  assign controls_horizontalDirectionValid = CICC1851_controls_frameStart[55];
  assign controls_verticalDirectionValid = CICC1851_controls_frameStart[56];
  assign controls_mainDirectionValid = CICC1851_controls_frameStart[57];
  assign controls_counterDirectionValid = CICC1851_controls_frameStart[58];
  assign controls_inValidMinDiff = CICC1851_controls_frameStart[59];
  always @(*) begin
    validStream_ready = (controlStream_ready && startRead);
    validStream_ready = (mainPixelAddrOneStream_ready && startRead);
    validStream_ready = (counterPixelAddrOneStream_ready && startRead);
    validStream_ready = (mainPixelAddrTwoStream_ready && startRead);
    validStream_ready = (counterPixelAddrTwoStream_ready && startRead);
    validStream_ready = (mainPixelAddrThreeStream_ready && startRead);
    validStream_ready = (counterPixelAddrThreeStream_ready && startRead);
    validStream_ready = (mainValidAddrOneStream_ready && startRead);
    validStream_ready = (counterValidAddrOneStream_ready && startRead);
    validStream_ready = (mainValidAddrTwoStream_ready && startRead);
    validStream_ready = (counterValidAddrTwoStream_ready && startRead);
    validStream_ready = (mainValidAddrThreeStream_ready && startRead);
    validStream_ready = (counterValidAddrThreeStream_ready && startRead);
  end

  assign controlStream_valid = (validStream_valid && startRead);
  assign controlStream_payload_frameStart = controls_frameStart;
  assign controlStream_payload_rowEnd = controls_rowEnd;
  assign controlStream_payload_pipeValid = controls_pipeValid;
  assign controlStream_payload_firstRow = controls_firstRow;
  assign controlStream_payload_lastRow = controls_lastRow;
  assign controlStream_payload_finalResult = controls_finalResult;
  assign controlStream_payload_mainCompare = controls_mainCompare;
  assign controlStream_payload_counterCompare = controls_counterCompare;
  assign controlStream_payload_horizontalCompare = controls_horizontalCompare;
  assign controlStream_payload_verticalCompare = controls_verticalCompare;
  assign controlStream_payload_mainDiff = controls_mainDiff;
  assign controlStream_payload_counterDiff = controls_counterDiff;
  assign controlStream_payload_horizontalDiff = controls_horizontalDiff;
  assign controlStream_payload_verticalDiff = controls_verticalDiff;
  assign controlStream_payload_isHorizontalMin = controls_isHorizontalMin;
  assign controlStream_payload_minDiff = controls_minDiff;
  assign controlStream_payload_currentPosition = controls_currentPosition;
  assign controlStream_payload_nextPosition = controls_nextPosition;
  assign controlStream_payload_horizontalDirectionValid = controls_horizontalDirectionValid;
  assign controlStream_payload_verticalDirectionValid = controls_verticalDirectionValid;
  assign controlStream_payload_mainDirectionValid = controls_mainDirectionValid;
  assign controlStream_payload_counterDirectionValid = controls_counterDirectionValid;
  assign controlStream_payload_inValidMinDiff = controls_inValidMinDiff;
  assign mainPixelAddrOneStream_valid = (validStream_valid && startRead);
  assign mainPixelAddrOneStream_payload = mainAddrOne;
  assign counterPixelAddrOneStream_valid = (validStream_valid && startRead);
  assign counterPixelAddrOneStream_payload = counterAddrOne;
  assign mainPixelAddrTwoStream_valid = (validStream_valid && startRead);
  assign mainPixelAddrTwoStream_payload = mainAddrTwo;
  assign counterPixelAddrTwoStream_valid = (validStream_valid && startRead);
  assign counterPixelAddrTwoStream_payload = counterAddrTwo;
  assign mainPixelAddrThreeStream_valid = (validStream_valid && startRead);
  assign mainPixelAddrThreeStream_payload = mainAddrThree;
  assign counterPixelAddrThreeStream_valid = (validStream_valid && startRead);
  assign counterPixelAddrThreeStream_payload = counterAddrThree;
  assign mainValidAddrOneStream_valid = (validStream_valid && startRead);
  assign mainValidAddrOneStream_payload = mainAddrOne;
  assign counterValidAddrOneStream_valid = (validStream_valid && startRead);
  assign counterValidAddrOneStream_payload = counterAddrOne;
  assign mainValidAddrTwoStream_valid = (validStream_valid && startRead);
  assign mainValidAddrTwoStream_payload = mainAddrTwo;
  assign counterValidAddrTwoStream_valid = (validStream_valid && startRead);
  assign counterValidAddrTwoStream_payload = counterAddrTwo;
  assign mainValidAddrThreeStream_valid = (validStream_valid && startRead);
  assign mainValidAddrThreeStream_payload = mainAddrThree;
  assign counterValidAddrThreeStream_valid = (validStream_valid && startRead);
  assign counterValidAddrThreeStream_payload = counterAddrThree;
  assign pixelsIn_s2mPipe_valid = (pixelsIn_valid || pixelsIn_rValid);
  assign pixelsIn_s2mPipe_payload_pixel = (pixelsIn_rValid ? pixelsIn_rData_pixel : pixelsIn_payload_pixel);
  assign pixelsIn_s2mPipe_payload_frameStart = (pixelsIn_rValid ? pixelsIn_rData_frameStart : pixelsIn_payload_frameStart);
  assign pixelsIn_s2mPipe_payload_rowEnd = (pixelsIn_rValid ? pixelsIn_rData_rowEnd : pixelsIn_payload_rowEnd);
  assign pixelsIn_s2mPipe_payload_inpValid = (pixelsIn_rValid ? pixelsIn_rData_inpValid : pixelsIn_payload_inpValid);
  always @(*) begin
    pixelsIn_s2mPipe_ready = pixelsIn_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368) begin
      pixelsIn_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368 = (! pixelsIn_s2mPipe_m2sPipe_valid);
  assign pixelsIn_s2mPipe_m2sPipe_valid = pixelsIn_s2mPipe_rValid;
  assign pixelsIn_s2mPipe_m2sPipe_payload_pixel = pixelsIn_s2mPipe_rData_pixel;
  assign pixelsIn_s2mPipe_m2sPipe_payload_frameStart = pixelsIn_s2mPipe_rData_frameStart;
  assign pixelsIn_s2mPipe_m2sPipe_payload_rowEnd = pixelsIn_s2mPipe_rData_rowEnd;
  assign pixelsIn_s2mPipe_m2sPipe_payload_inpValid = pixelsIn_s2mPipe_rData_inpValid;
  assign passPixels_valid = (pixelsIn_s2mPipe_m2sPipe_valid && bufferEnable);
  assign pixelsIn_s2mPipe_m2sPipe_ready = (passPixels_ready && bufferEnable);
  assign passPixels_payload_pixel = pixelsIn_s2mPipe_m2sPipe_payload_pixel;
  assign passPixels_payload_frameStart = pixelsIn_s2mPipe_m2sPipe_payload_frameStart;
  assign passPixels_payload_rowEnd = pixelsIn_s2mPipe_m2sPipe_payload_rowEnd;
  assign passPixels_payload_inpValid = pixelsIn_s2mPipe_m2sPipe_payload_inpValid;
  assign passPixels_ready = 1'b1;
  assign passPixels_fire = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart3_l226 = ((CICC1851_when_SuperResolutionPart3_l226 == CICC1851_when_SuperResolutionPart3_l226_1) && passPixels_fire);
  assign passPixels_fire_1 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart3_l227 = (((CICC1851_when_SuperResolutionPart3_l227 == CICC1851_when_SuperResolutionPart3_l227_1) && bufferReachRowEnd) && passPixels_fire_1);
  assign passPixels_fire_2 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart3_l230 = (passPixels_payload_rowEnd && passPixels_fire_2);
  assign passPixels_fire_3 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart3_l243 = (passPixels_payload_rowEnd && passPixels_fire_3);
  assign when_SuperResolutionPart3_l244 = (bufferSwitch == 2'b10);
  assign passPixels_fire_4 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart3_l251 = (((12'h002 <= bufferRowCount_value) && passPixels_payload_rowEnd) && passPixels_fire_4);
  assign when_SuperResolutionPart3_l255 = (bufferReachFinalRow && bufferReachRowEnd);
  assign passPixels_fire_5 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart3_l262 = (passPixels_payload_frameStart && passPixels_fire_5);
  assign pixelsOut_fire = (pixelsOut_valid && pixelsOut_ready);
  assign when_SuperResolutionPart3_l270 = ((CICC1851_when_SuperResolutionPart3_l270 == CICC1851_when_SuperResolutionPart3_l270_1) && pixelsOut_fire);
  assign pixelsOut_fire_1 = (pixelsOut_valid && pixelsOut_ready);
  assign when_SuperResolutionPart3_l271 = (((CICC1851_when_SuperResolutionPart3_l271 == CICC1851_when_SuperResolutionPart3_l271_1) && alreadyReachRowEnd) && pixelsOut_fire_1);
  assign pixelsOut_fire_2 = (pixelsOut_valid && pixelsOut_ready);
  assign pixelsOut_fire_3 = (pixelsOut_valid && pixelsOut_ready);
  assign when_SuperResolutionPart3_l282 = ((alreadyReachFinalRow && alreadyReachRowEnd) && pixelsOut_fire_3);
  assign passPixels_fire_6 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_7 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_8 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_9 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_10 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_11 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_12 = (passPixels_valid && passPixels_ready);
  assign mainPixelAddrOneStream_ready = (! mainPixelAddrOneStream_rValid);
  assign mainPixelAddrOneStream_s2mPipe_valid = (mainPixelAddrOneStream_valid || mainPixelAddrOneStream_rValid);
  assign mainPixelAddrOneStream_s2mPipe_payload = (mainPixelAddrOneStream_rValid ? mainPixelAddrOneStream_rData : mainPixelAddrOneStream_payload);
  always @(*) begin
    mainPixelAddrOneStream_s2mPipe_ready = mainPixelAddrOneStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_1) begin
      mainPixelAddrOneStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_1 = (! mainPixelAddrOneStream_s2mPipe_m2sPipe_valid);
  assign mainPixelAddrOneStream_s2mPipe_m2sPipe_valid = mainPixelAddrOneStream_s2mPipe_rValid;
  assign mainPixelAddrOneStream_s2mPipe_m2sPipe_payload = mainPixelAddrOneStream_s2mPipe_rData;
  assign mainPixelAddrOneStream_s2mPipe_m2sPipe_ready = ((! CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready) || CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready = CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_mainOnePixelStream_payload = CICC1851_lineBufferOne_port1;
  assign CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_1 = readStage_mainOnePixelStream_ready;
    if(when_Stream_l368_2) begin
      CICC1851_1 = 1'b1;
    end
  end

  assign when_Stream_l368_2 = (! readStage_mainOnePixelStream_valid);
  assign readStage_mainOnePixelStream_valid = CICC1851_readStage_mainOnePixelStream_valid;
  assign readStage_mainOnePixelStream_payload = CICC1851_readStage_mainOnePixelStream_payload_2;
  assign counterPixelAddrOneStream_ready = (! counterPixelAddrOneStream_rValid);
  assign counterPixelAddrOneStream_s2mPipe_valid = (counterPixelAddrOneStream_valid || counterPixelAddrOneStream_rValid);
  assign counterPixelAddrOneStream_s2mPipe_payload = (counterPixelAddrOneStream_rValid ? counterPixelAddrOneStream_rData : counterPixelAddrOneStream_payload);
  always @(*) begin
    counterPixelAddrOneStream_s2mPipe_ready = counterPixelAddrOneStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_3) begin
      counterPixelAddrOneStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_3 = (! counterPixelAddrOneStream_s2mPipe_m2sPipe_valid);
  assign counterPixelAddrOneStream_s2mPipe_m2sPipe_valid = counterPixelAddrOneStream_s2mPipe_rValid;
  assign counterPixelAddrOneStream_s2mPipe_m2sPipe_payload = counterPixelAddrOneStream_s2mPipe_rData;
  assign counterPixelAddrOneStream_s2mPipe_m2sPipe_ready = ((! CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready) || CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready = CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_counterOnePixelStream_payload = CICC1851_lineBufferOne_port2;
  assign CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_2 = readStage_counterOnePixelStream_ready;
    if(when_Stream_l368_4) begin
      CICC1851_2 = 1'b1;
    end
  end

  assign when_Stream_l368_4 = (! readStage_counterOnePixelStream_valid);
  assign readStage_counterOnePixelStream_valid = CICC1851_readStage_counterOnePixelStream_valid;
  assign readStage_counterOnePixelStream_payload = CICC1851_readStage_counterOnePixelStream_payload_2;
  assign mainPixelAddrTwoStream_ready = (! mainPixelAddrTwoStream_rValid);
  assign mainPixelAddrTwoStream_s2mPipe_valid = (mainPixelAddrTwoStream_valid || mainPixelAddrTwoStream_rValid);
  assign mainPixelAddrTwoStream_s2mPipe_payload = (mainPixelAddrTwoStream_rValid ? mainPixelAddrTwoStream_rData : mainPixelAddrTwoStream_payload);
  always @(*) begin
    mainPixelAddrTwoStream_s2mPipe_ready = mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_5) begin
      mainPixelAddrTwoStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_5 = (! mainPixelAddrTwoStream_s2mPipe_m2sPipe_valid);
  assign mainPixelAddrTwoStream_s2mPipe_m2sPipe_valid = mainPixelAddrTwoStream_s2mPipe_rValid;
  assign mainPixelAddrTwoStream_s2mPipe_m2sPipe_payload = mainPixelAddrTwoStream_s2mPipe_rData;
  assign mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready = ((! CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready) || CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready = CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_mainTwoPixelStream_payload = CICC1851_lineBufferTwo_port1;
  assign CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_3 = readStage_mainTwoPixelStream_ready;
    if(when_Stream_l368_6) begin
      CICC1851_3 = 1'b1;
    end
  end

  assign when_Stream_l368_6 = (! readStage_mainTwoPixelStream_valid);
  assign readStage_mainTwoPixelStream_valid = CICC1851_readStage_mainTwoPixelStream_valid;
  assign readStage_mainTwoPixelStream_payload = CICC1851_readStage_mainTwoPixelStream_payload_2;
  assign counterPixelAddrTwoStream_ready = (! counterPixelAddrTwoStream_rValid);
  assign counterPixelAddrTwoStream_s2mPipe_valid = (counterPixelAddrTwoStream_valid || counterPixelAddrTwoStream_rValid);
  assign counterPixelAddrTwoStream_s2mPipe_payload = (counterPixelAddrTwoStream_rValid ? counterPixelAddrTwoStream_rData : counterPixelAddrTwoStream_payload);
  always @(*) begin
    counterPixelAddrTwoStream_s2mPipe_ready = counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_7) begin
      counterPixelAddrTwoStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_7 = (! counterPixelAddrTwoStream_s2mPipe_m2sPipe_valid);
  assign counterPixelAddrTwoStream_s2mPipe_m2sPipe_valid = counterPixelAddrTwoStream_s2mPipe_rValid;
  assign counterPixelAddrTwoStream_s2mPipe_m2sPipe_payload = counterPixelAddrTwoStream_s2mPipe_rData;
  assign counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready = ((! CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready) || CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready = CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_counterTwoPixelStream_payload = CICC1851_lineBufferTwo_port2;
  assign CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_4 = readStage_counterTwoPixelStream_ready;
    if(when_Stream_l368_8) begin
      CICC1851_4 = 1'b1;
    end
  end

  assign when_Stream_l368_8 = (! readStage_counterTwoPixelStream_valid);
  assign readStage_counterTwoPixelStream_valid = CICC1851_readStage_counterTwoPixelStream_valid;
  assign readStage_counterTwoPixelStream_payload = CICC1851_readStage_counterTwoPixelStream_payload_2;
  assign mainPixelAddrThreeStream_ready = (! mainPixelAddrThreeStream_rValid);
  assign mainPixelAddrThreeStream_s2mPipe_valid = (mainPixelAddrThreeStream_valid || mainPixelAddrThreeStream_rValid);
  assign mainPixelAddrThreeStream_s2mPipe_payload = (mainPixelAddrThreeStream_rValid ? mainPixelAddrThreeStream_rData : mainPixelAddrThreeStream_payload);
  always @(*) begin
    mainPixelAddrThreeStream_s2mPipe_ready = mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_9) begin
      mainPixelAddrThreeStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_9 = (! mainPixelAddrThreeStream_s2mPipe_m2sPipe_valid);
  assign mainPixelAddrThreeStream_s2mPipe_m2sPipe_valid = mainPixelAddrThreeStream_s2mPipe_rValid;
  assign mainPixelAddrThreeStream_s2mPipe_m2sPipe_payload = mainPixelAddrThreeStream_s2mPipe_rData;
  assign mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready = ((! CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready) || CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready = CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_mainThreePixelStream_payload = CICC1851_lineBufferThree_port1;
  assign CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_5 = readStage_mainThreePixelStream_ready;
    if(when_Stream_l368_10) begin
      CICC1851_5 = 1'b1;
    end
  end

  assign when_Stream_l368_10 = (! readStage_mainThreePixelStream_valid);
  assign readStage_mainThreePixelStream_valid = CICC1851_readStage_mainThreePixelStream_valid;
  assign readStage_mainThreePixelStream_payload = CICC1851_readStage_mainThreePixelStream_payload_2;
  assign counterPixelAddrThreeStream_ready = (! counterPixelAddrThreeStream_rValid);
  assign counterPixelAddrThreeStream_s2mPipe_valid = (counterPixelAddrThreeStream_valid || counterPixelAddrThreeStream_rValid);
  assign counterPixelAddrThreeStream_s2mPipe_payload = (counterPixelAddrThreeStream_rValid ? counterPixelAddrThreeStream_rData : counterPixelAddrThreeStream_payload);
  always @(*) begin
    counterPixelAddrThreeStream_s2mPipe_ready = counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_11) begin
      counterPixelAddrThreeStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_11 = (! counterPixelAddrThreeStream_s2mPipe_m2sPipe_valid);
  assign counterPixelAddrThreeStream_s2mPipe_m2sPipe_valid = counterPixelAddrThreeStream_s2mPipe_rValid;
  assign counterPixelAddrThreeStream_s2mPipe_m2sPipe_payload = counterPixelAddrThreeStream_s2mPipe_rData;
  assign counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready = ((! CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready) || CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready = CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_counterThreePixelStream_payload = CICC1851_lineBufferThree_port2;
  assign CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_6 = readStage_counterThreePixelStream_ready;
    if(when_Stream_l368_12) begin
      CICC1851_6 = 1'b1;
    end
  end

  assign when_Stream_l368_12 = (! readStage_counterThreePixelStream_valid);
  assign readStage_counterThreePixelStream_valid = CICC1851_readStage_counterThreePixelStream_valid;
  assign readStage_counterThreePixelStream_payload = CICC1851_readStage_counterThreePixelStream_payload_2;
  assign mainValidAddrOneStream_ready = (! mainValidAddrOneStream_rValid);
  assign mainValidAddrOneStream_s2mPipe_valid = (mainValidAddrOneStream_valid || mainValidAddrOneStream_rValid);
  assign mainValidAddrOneStream_s2mPipe_payload = (mainValidAddrOneStream_rValid ? mainValidAddrOneStream_rData : mainValidAddrOneStream_payload);
  always @(*) begin
    mainValidAddrOneStream_s2mPipe_ready = mainValidAddrOneStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_13) begin
      mainValidAddrOneStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_13 = (! mainValidAddrOneStream_s2mPipe_m2sPipe_valid);
  assign mainValidAddrOneStream_s2mPipe_m2sPipe_valid = mainValidAddrOneStream_s2mPipe_rValid;
  assign mainValidAddrOneStream_s2mPipe_m2sPipe_payload = mainValidAddrOneStream_s2mPipe_rData;
  assign mainValidAddrOneStream_s2mPipe_m2sPipe_ready = ((! CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready) || CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready = CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_mainOneValidStream_payload = CICC1851_validBufferOne_port1[0];
  assign CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_7 = readStage_mainOneValidStream_ready;
    if(when_Stream_l368_14) begin
      CICC1851_7 = 1'b1;
    end
  end

  assign when_Stream_l368_14 = (! readStage_mainOneValidStream_valid);
  assign readStage_mainOneValidStream_valid = CICC1851_readStage_mainOneValidStream_valid;
  assign readStage_mainOneValidStream_payload = CICC1851_readStage_mainOneValidStream_payload_2;
  assign counterValidAddrOneStream_ready = (! counterValidAddrOneStream_rValid);
  assign counterValidAddrOneStream_s2mPipe_valid = (counterValidAddrOneStream_valid || counterValidAddrOneStream_rValid);
  assign counterValidAddrOneStream_s2mPipe_payload = (counterValidAddrOneStream_rValid ? counterValidAddrOneStream_rData : counterValidAddrOneStream_payload);
  always @(*) begin
    counterValidAddrOneStream_s2mPipe_ready = counterValidAddrOneStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_15) begin
      counterValidAddrOneStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_15 = (! counterValidAddrOneStream_s2mPipe_m2sPipe_valid);
  assign counterValidAddrOneStream_s2mPipe_m2sPipe_valid = counterValidAddrOneStream_s2mPipe_rValid;
  assign counterValidAddrOneStream_s2mPipe_m2sPipe_payload = counterValidAddrOneStream_s2mPipe_rData;
  assign counterValidAddrOneStream_s2mPipe_m2sPipe_ready = ((! CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready) || CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready = CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_counterOneValidStream_payload = CICC1851_validBufferOne_port2[0];
  assign CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_8 = readStage_counterOneValidStream_ready;
    if(when_Stream_l368_16) begin
      CICC1851_8 = 1'b1;
    end
  end

  assign when_Stream_l368_16 = (! readStage_counterOneValidStream_valid);
  assign readStage_counterOneValidStream_valid = CICC1851_readStage_counterOneValidStream_valid;
  assign readStage_counterOneValidStream_payload = CICC1851_readStage_counterOneValidStream_payload_2;
  assign mainValidAddrTwoStream_ready = (! mainValidAddrTwoStream_rValid);
  assign mainValidAddrTwoStream_s2mPipe_valid = (mainValidAddrTwoStream_valid || mainValidAddrTwoStream_rValid);
  assign mainValidAddrTwoStream_s2mPipe_payload = (mainValidAddrTwoStream_rValid ? mainValidAddrTwoStream_rData : mainValidAddrTwoStream_payload);
  always @(*) begin
    mainValidAddrTwoStream_s2mPipe_ready = mainValidAddrTwoStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_17) begin
      mainValidAddrTwoStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_17 = (! mainValidAddrTwoStream_s2mPipe_m2sPipe_valid);
  assign mainValidAddrTwoStream_s2mPipe_m2sPipe_valid = mainValidAddrTwoStream_s2mPipe_rValid;
  assign mainValidAddrTwoStream_s2mPipe_m2sPipe_payload = mainValidAddrTwoStream_s2mPipe_rData;
  assign mainValidAddrTwoStream_s2mPipe_m2sPipe_ready = ((! CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready) || CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready = CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_mainTwoValidStream_payload = CICC1851_validBufferTwo_port1[0];
  assign CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_9 = readStage_mainTwoValidStream_ready;
    if(when_Stream_l368_18) begin
      CICC1851_9 = 1'b1;
    end
  end

  assign when_Stream_l368_18 = (! readStage_mainTwoValidStream_valid);
  assign readStage_mainTwoValidStream_valid = CICC1851_readStage_mainTwoValidStream_valid;
  assign readStage_mainTwoValidStream_payload = CICC1851_readStage_mainTwoValidStream_payload_2;
  assign counterValidAddrTwoStream_ready = (! counterValidAddrTwoStream_rValid);
  assign counterValidAddrTwoStream_s2mPipe_valid = (counterValidAddrTwoStream_valid || counterValidAddrTwoStream_rValid);
  assign counterValidAddrTwoStream_s2mPipe_payload = (counterValidAddrTwoStream_rValid ? counterValidAddrTwoStream_rData : counterValidAddrTwoStream_payload);
  always @(*) begin
    counterValidAddrTwoStream_s2mPipe_ready = counterValidAddrTwoStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_19) begin
      counterValidAddrTwoStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_19 = (! counterValidAddrTwoStream_s2mPipe_m2sPipe_valid);
  assign counterValidAddrTwoStream_s2mPipe_m2sPipe_valid = counterValidAddrTwoStream_s2mPipe_rValid;
  assign counterValidAddrTwoStream_s2mPipe_m2sPipe_payload = counterValidAddrTwoStream_s2mPipe_rData;
  assign counterValidAddrTwoStream_s2mPipe_m2sPipe_ready = ((! CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready) || CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready = CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_counterTwoValidStream_payload = CICC1851_validBufferTwo_port2[0];
  assign CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_10 = readStage_counterTwoValidStream_ready;
    if(when_Stream_l368_20) begin
      CICC1851_10 = 1'b1;
    end
  end

  assign when_Stream_l368_20 = (! readStage_counterTwoValidStream_valid);
  assign readStage_counterTwoValidStream_valid = CICC1851_readStage_counterTwoValidStream_valid;
  assign readStage_counterTwoValidStream_payload = CICC1851_readStage_counterTwoValidStream_payload_2;
  assign mainValidAddrThreeStream_ready = (! mainValidAddrThreeStream_rValid);
  assign mainValidAddrThreeStream_s2mPipe_valid = (mainValidAddrThreeStream_valid || mainValidAddrThreeStream_rValid);
  assign mainValidAddrThreeStream_s2mPipe_payload = (mainValidAddrThreeStream_rValid ? mainValidAddrThreeStream_rData : mainValidAddrThreeStream_payload);
  always @(*) begin
    mainValidAddrThreeStream_s2mPipe_ready = mainValidAddrThreeStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_21) begin
      mainValidAddrThreeStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_21 = (! mainValidAddrThreeStream_s2mPipe_m2sPipe_valid);
  assign mainValidAddrThreeStream_s2mPipe_m2sPipe_valid = mainValidAddrThreeStream_s2mPipe_rValid;
  assign mainValidAddrThreeStream_s2mPipe_m2sPipe_payload = mainValidAddrThreeStream_s2mPipe_rData;
  assign mainValidAddrThreeStream_s2mPipe_m2sPipe_ready = ((! CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready) || CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready = CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_mainThreeValidStream_payload = CICC1851_validBufferThree_port1[0];
  assign CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_11 = readStage_mainThreeValidStream_ready;
    if(when_Stream_l368_22) begin
      CICC1851_11 = 1'b1;
    end
  end

  assign when_Stream_l368_22 = (! readStage_mainThreeValidStream_valid);
  assign readStage_mainThreeValidStream_valid = CICC1851_readStage_mainThreeValidStream_valid;
  assign readStage_mainThreeValidStream_payload = CICC1851_readStage_mainThreeValidStream_payload_2;
  assign counterValidAddrThreeStream_ready = (! counterValidAddrThreeStream_rValid);
  assign counterValidAddrThreeStream_s2mPipe_valid = (counterValidAddrThreeStream_valid || counterValidAddrThreeStream_rValid);
  assign counterValidAddrThreeStream_s2mPipe_payload = (counterValidAddrThreeStream_rValid ? counterValidAddrThreeStream_rData : counterValidAddrThreeStream_payload);
  always @(*) begin
    counterValidAddrThreeStream_s2mPipe_ready = counterValidAddrThreeStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_23) begin
      counterValidAddrThreeStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_23 = (! counterValidAddrThreeStream_s2mPipe_m2sPipe_valid);
  assign counterValidAddrThreeStream_s2mPipe_m2sPipe_valid = counterValidAddrThreeStream_s2mPipe_rValid;
  assign counterValidAddrThreeStream_s2mPipe_m2sPipe_payload = counterValidAddrThreeStream_s2mPipe_rData;
  assign counterValidAddrThreeStream_s2mPipe_m2sPipe_ready = ((! CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready) || CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready = CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_counterThreeValidStream_payload = CICC1851_validBufferThree_port2[0];
  assign CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_12 = readStage_counterThreeValidStream_ready;
    if(when_Stream_l368_24) begin
      CICC1851_12 = 1'b1;
    end
  end

  assign when_Stream_l368_24 = (! readStage_counterThreeValidStream_valid);
  assign readStage_counterThreeValidStream_valid = CICC1851_readStage_counterThreeValidStream_valid;
  assign readStage_counterThreeValidStream_payload = CICC1851_readStage_counterThreeValidStream_payload_2;
  assign controlStream_ready = (! controlStream_rValid);
  assign controlStream_s2mPipe_valid = (controlStream_valid || controlStream_rValid);
  assign controlStream_s2mPipe_payload_frameStart = (controlStream_rValid ? controlStream_rData_frameStart : controlStream_payload_frameStart);
  assign controlStream_s2mPipe_payload_rowEnd = (controlStream_rValid ? controlStream_rData_rowEnd : controlStream_payload_rowEnd);
  assign controlStream_s2mPipe_payload_pipeValid = (controlStream_rValid ? controlStream_rData_pipeValid : controlStream_payload_pipeValid);
  assign controlStream_s2mPipe_payload_firstRow = (controlStream_rValid ? controlStream_rData_firstRow : controlStream_payload_firstRow);
  assign controlStream_s2mPipe_payload_lastRow = (controlStream_rValid ? controlStream_rData_lastRow : controlStream_payload_lastRow);
  assign controlStream_s2mPipe_payload_finalResult = (controlStream_rValid ? controlStream_rData_finalResult : controlStream_payload_finalResult);
  assign controlStream_s2mPipe_payload_mainCompare = (controlStream_rValid ? controlStream_rData_mainCompare : controlStream_payload_mainCompare);
  assign controlStream_s2mPipe_payload_counterCompare = (controlStream_rValid ? controlStream_rData_counterCompare : controlStream_payload_counterCompare);
  assign controlStream_s2mPipe_payload_horizontalCompare = (controlStream_rValid ? controlStream_rData_horizontalCompare : controlStream_payload_horizontalCompare);
  assign controlStream_s2mPipe_payload_verticalCompare = (controlStream_rValid ? controlStream_rData_verticalCompare : controlStream_payload_verticalCompare);
  assign controlStream_s2mPipe_payload_mainDiff = (controlStream_rValid ? controlStream_rData_mainDiff : controlStream_payload_mainDiff);
  assign controlStream_s2mPipe_payload_counterDiff = (controlStream_rValid ? controlStream_rData_counterDiff : controlStream_payload_counterDiff);
  assign controlStream_s2mPipe_payload_horizontalDiff = (controlStream_rValid ? controlStream_rData_horizontalDiff : controlStream_payload_horizontalDiff);
  assign controlStream_s2mPipe_payload_verticalDiff = (controlStream_rValid ? controlStream_rData_verticalDiff : controlStream_payload_verticalDiff);
  assign controlStream_s2mPipe_payload_isHorizontalMin = (controlStream_rValid ? controlStream_rData_isHorizontalMin : controlStream_payload_isHorizontalMin);
  assign controlStream_s2mPipe_payload_minDiff = (controlStream_rValid ? controlStream_rData_minDiff : controlStream_payload_minDiff);
  assign controlStream_s2mPipe_payload_currentPosition = (controlStream_rValid ? controlStream_rData_currentPosition : controlStream_payload_currentPosition);
  assign controlStream_s2mPipe_payload_nextPosition = (controlStream_rValid ? controlStream_rData_nextPosition : controlStream_payload_nextPosition);
  assign controlStream_s2mPipe_payload_horizontalDirectionValid = (controlStream_rValid ? controlStream_rData_horizontalDirectionValid : controlStream_payload_horizontalDirectionValid);
  assign controlStream_s2mPipe_payload_verticalDirectionValid = (controlStream_rValid ? controlStream_rData_verticalDirectionValid : controlStream_payload_verticalDirectionValid);
  assign controlStream_s2mPipe_payload_mainDirectionValid = (controlStream_rValid ? controlStream_rData_mainDirectionValid : controlStream_payload_mainDirectionValid);
  assign controlStream_s2mPipe_payload_counterDirectionValid = (controlStream_rValid ? controlStream_rData_counterDirectionValid : controlStream_payload_counterDirectionValid);
  assign controlStream_s2mPipe_payload_inValidMinDiff = (controlStream_rValid ? controlStream_rData_inValidMinDiff : controlStream_payload_inValidMinDiff);
  always @(*) begin
    controlStream_s2mPipe_ready = controlStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_25) begin
      controlStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_25 = (! controlStream_s2mPipe_m2sPipe_valid);
  assign controlStream_s2mPipe_m2sPipe_valid = controlStream_s2mPipe_rValid;
  assign controlStream_s2mPipe_m2sPipe_payload_frameStart = controlStream_s2mPipe_rData_frameStart;
  assign controlStream_s2mPipe_m2sPipe_payload_rowEnd = controlStream_s2mPipe_rData_rowEnd;
  assign controlStream_s2mPipe_m2sPipe_payload_pipeValid = controlStream_s2mPipe_rData_pipeValid;
  assign controlStream_s2mPipe_m2sPipe_payload_firstRow = controlStream_s2mPipe_rData_firstRow;
  assign controlStream_s2mPipe_m2sPipe_payload_lastRow = controlStream_s2mPipe_rData_lastRow;
  assign controlStream_s2mPipe_m2sPipe_payload_finalResult = controlStream_s2mPipe_rData_finalResult;
  assign controlStream_s2mPipe_m2sPipe_payload_mainCompare = controlStream_s2mPipe_rData_mainCompare;
  assign controlStream_s2mPipe_m2sPipe_payload_counterCompare = controlStream_s2mPipe_rData_counterCompare;
  assign controlStream_s2mPipe_m2sPipe_payload_horizontalCompare = controlStream_s2mPipe_rData_horizontalCompare;
  assign controlStream_s2mPipe_m2sPipe_payload_verticalCompare = controlStream_s2mPipe_rData_verticalCompare;
  assign controlStream_s2mPipe_m2sPipe_payload_mainDiff = controlStream_s2mPipe_rData_mainDiff;
  assign controlStream_s2mPipe_m2sPipe_payload_counterDiff = controlStream_s2mPipe_rData_counterDiff;
  assign controlStream_s2mPipe_m2sPipe_payload_horizontalDiff = controlStream_s2mPipe_rData_horizontalDiff;
  assign controlStream_s2mPipe_m2sPipe_payload_verticalDiff = controlStream_s2mPipe_rData_verticalDiff;
  assign controlStream_s2mPipe_m2sPipe_payload_isHorizontalMin = controlStream_s2mPipe_rData_isHorizontalMin;
  assign controlStream_s2mPipe_m2sPipe_payload_minDiff = controlStream_s2mPipe_rData_minDiff;
  assign controlStream_s2mPipe_m2sPipe_payload_currentPosition = controlStream_s2mPipe_rData_currentPosition;
  assign controlStream_s2mPipe_m2sPipe_payload_nextPosition = controlStream_s2mPipe_rData_nextPosition;
  assign controlStream_s2mPipe_m2sPipe_payload_horizontalDirectionValid = controlStream_s2mPipe_rData_horizontalDirectionValid;
  assign controlStream_s2mPipe_m2sPipe_payload_verticalDirectionValid = controlStream_s2mPipe_rData_verticalDirectionValid;
  assign controlStream_s2mPipe_m2sPipe_payload_mainDirectionValid = controlStream_s2mPipe_rData_mainDirectionValid;
  assign controlStream_s2mPipe_m2sPipe_payload_counterDirectionValid = controlStream_s2mPipe_rData_counterDirectionValid;
  assign controlStream_s2mPipe_m2sPipe_payload_inValidMinDiff = controlStream_s2mPipe_rData_inValidMinDiff;
  always @(*) begin
    controlStream_s2mPipe_m2sPipe_ready = controlStream_s2mPipe_m2sPipe_m2sPipe_ready;
    if(when_Stream_l368_26) begin
      controlStream_s2mPipe_m2sPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_26 = (! controlStream_s2mPipe_m2sPipe_m2sPipe_valid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_valid = controlStream_s2mPipe_m2sPipe_rValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_frameStart = controlStream_s2mPipe_m2sPipe_rData_frameStart;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_rowEnd = controlStream_s2mPipe_m2sPipe_rData_rowEnd;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_pipeValid = controlStream_s2mPipe_m2sPipe_rData_pipeValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_firstRow = controlStream_s2mPipe_m2sPipe_rData_firstRow;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_lastRow = controlStream_s2mPipe_m2sPipe_rData_lastRow;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_finalResult = controlStream_s2mPipe_m2sPipe_rData_finalResult;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainCompare = controlStream_s2mPipe_m2sPipe_rData_mainCompare;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterCompare = controlStream_s2mPipe_m2sPipe_rData_counterCompare;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_horizontalCompare = controlStream_s2mPipe_m2sPipe_rData_horizontalCompare;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_verticalCompare = controlStream_s2mPipe_m2sPipe_rData_verticalCompare;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDiff = controlStream_s2mPipe_m2sPipe_rData_mainDiff;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDiff = controlStream_s2mPipe_m2sPipe_rData_counterDiff;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_horizontalDiff = controlStream_s2mPipe_m2sPipe_rData_horizontalDiff;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_verticalDiff = controlStream_s2mPipe_m2sPipe_rData_verticalDiff;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_isHorizontalMin = controlStream_s2mPipe_m2sPipe_rData_isHorizontalMin;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_minDiff = controlStream_s2mPipe_m2sPipe_rData_minDiff;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_currentPosition = controlStream_s2mPipe_m2sPipe_rData_currentPosition;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_nextPosition = controlStream_s2mPipe_m2sPipe_rData_nextPosition;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_horizontalDirectionValid = controlStream_s2mPipe_m2sPipe_rData_horizontalDirectionValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_verticalDirectionValid = controlStream_s2mPipe_m2sPipe_rData_verticalDirectionValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDirectionValid = controlStream_s2mPipe_m2sPipe_rData_mainDirectionValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDirectionValid = controlStream_s2mPipe_m2sPipe_rData_counterDirectionValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_inValidMinDiff = controlStream_s2mPipe_m2sPipe_rData_inValidMinDiff;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_ready = (! controlStream_s2mPipe_m2sPipe_m2sPipe_rValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_valid = (controlStream_s2mPipe_m2sPipe_m2sPipe_valid || controlStream_s2mPipe_m2sPipe_m2sPipe_rValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_frameStart = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_frameStart : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_frameStart);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_rowEnd = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_rowEnd : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_rowEnd);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_pipeValid = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_pipeValid : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_pipeValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_firstRow = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_firstRow : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_firstRow);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_lastRow = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_lastRow : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_lastRow);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_finalResult = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_finalResult : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_finalResult);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainCompare = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainCompare : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainCompare);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterCompare = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterCompare : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterCompare);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_horizontalCompare = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_horizontalCompare : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_horizontalCompare);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_verticalCompare = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_verticalCompare : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_verticalCompare);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainDiff = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainDiff : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDiff);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterDiff = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterDiff : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDiff);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_horizontalDiff = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_horizontalDiff : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_horizontalDiff);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_verticalDiff = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_verticalDiff : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_verticalDiff);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_isHorizontalMin = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_isHorizontalMin : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_isHorizontalMin);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_minDiff = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_minDiff : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_minDiff);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_currentPosition = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_currentPosition : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_currentPosition);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_nextPosition = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_nextPosition : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_nextPosition);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_horizontalDirectionValid = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_horizontalDirectionValid : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_horizontalDirectionValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_verticalDirectionValid = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_verticalDirectionValid : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_verticalDirectionValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainDirectionValid = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainDirectionValid : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDirectionValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterDirectionValid = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterDirectionValid : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDirectionValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_inValidMinDiff = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_inValidMinDiff : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_inValidMinDiff);
  always @(*) begin
    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready = readStage_controlPipe_ready;
    if(when_Stream_l368_27) begin
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_27 = (! readStage_controlPipe_valid);
  assign readStage_controlPipe_valid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rValid;
  assign readStage_controlPipe_payload_frameStart = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_frameStart;
  assign readStage_controlPipe_payload_rowEnd = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_rowEnd;
  assign readStage_controlPipe_payload_pipeValid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_pipeValid;
  assign readStage_controlPipe_payload_firstRow = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_firstRow;
  assign readStage_controlPipe_payload_lastRow = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_lastRow;
  assign readStage_controlPipe_payload_finalResult = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_finalResult;
  assign readStage_controlPipe_payload_mainCompare = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainCompare;
  assign readStage_controlPipe_payload_counterCompare = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterCompare;
  assign readStage_controlPipe_payload_horizontalCompare = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_horizontalCompare;
  assign readStage_controlPipe_payload_verticalCompare = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_verticalCompare;
  assign readStage_controlPipe_payload_mainDiff = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainDiff;
  assign readStage_controlPipe_payload_counterDiff = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterDiff;
  assign readStage_controlPipe_payload_horizontalDiff = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_horizontalDiff;
  assign readStage_controlPipe_payload_verticalDiff = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_verticalDiff;
  assign readStage_controlPipe_payload_isHorizontalMin = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_isHorizontalMin;
  assign readStage_controlPipe_payload_minDiff = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_minDiff;
  assign readStage_controlPipe_payload_currentPosition = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_currentPosition;
  assign readStage_controlPipe_payload_nextPosition = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_nextPosition;
  assign readStage_controlPipe_payload_horizontalDirectionValid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_horizontalDirectionValid;
  assign readStage_controlPipe_payload_verticalDirectionValid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_verticalDirectionValid;
  assign readStage_controlPipe_payload_mainDirectionValid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainDirectionValid;
  assign readStage_controlPipe_payload_counterDirectionValid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterDirectionValid;
  assign readStage_controlPipe_payload_inValidMinDiff = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_inValidMinDiff;
  assign readStage_mainOnePixelStream_ready = (! readStage_mainOnePixelStream_rValid);
  assign readStage_mainOnePixelStream_s2mPipe_valid = (readStage_mainOnePixelStream_valid || readStage_mainOnePixelStream_rValid);
  assign readStage_mainOnePixelStream_s2mPipe_payload = (readStage_mainOnePixelStream_rValid ? readStage_mainOnePixelStream_rData : readStage_mainOnePixelStream_payload);
  always @(*) begin
    readStage_mainOnePixelStream_s2mPipe_ready = compareStage_mainOnePixelStream_ready;
    if(when_Stream_l368_28) begin
      readStage_mainOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_28 = (! compareStage_mainOnePixelStream_valid);
  assign compareStage_mainOnePixelStream_valid = readStage_mainOnePixelStream_s2mPipe_rValid;
  assign compareStage_mainOnePixelStream_payload = readStage_mainOnePixelStream_s2mPipe_rData;
  assign readStage_counterOnePixelStream_ready = (! readStage_counterOnePixelStream_rValid);
  assign readStage_counterOnePixelStream_s2mPipe_valid = (readStage_counterOnePixelStream_valid || readStage_counterOnePixelStream_rValid);
  assign readStage_counterOnePixelStream_s2mPipe_payload = (readStage_counterOnePixelStream_rValid ? readStage_counterOnePixelStream_rData : readStage_counterOnePixelStream_payload);
  always @(*) begin
    readStage_counterOnePixelStream_s2mPipe_ready = compareStage_counterOnePixelStream_ready;
    if(when_Stream_l368_29) begin
      readStage_counterOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_29 = (! compareStage_counterOnePixelStream_valid);
  assign compareStage_counterOnePixelStream_valid = readStage_counterOnePixelStream_s2mPipe_rValid;
  assign compareStage_counterOnePixelStream_payload = readStage_counterOnePixelStream_s2mPipe_rData;
  assign readStage_mainTwoPixelStream_ready = (! readStage_mainTwoPixelStream_rValid);
  assign readStage_mainTwoPixelStream_s2mPipe_valid = (readStage_mainTwoPixelStream_valid || readStage_mainTwoPixelStream_rValid);
  assign readStage_mainTwoPixelStream_s2mPipe_payload = (readStage_mainTwoPixelStream_rValid ? readStage_mainTwoPixelStream_rData : readStage_mainTwoPixelStream_payload);
  always @(*) begin
    readStage_mainTwoPixelStream_s2mPipe_ready = compareStage_mainTwoPixelStream_ready;
    if(when_Stream_l368_30) begin
      readStage_mainTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_30 = (! compareStage_mainTwoPixelStream_valid);
  assign compareStage_mainTwoPixelStream_valid = readStage_mainTwoPixelStream_s2mPipe_rValid;
  assign compareStage_mainTwoPixelStream_payload = readStage_mainTwoPixelStream_s2mPipe_rData;
  assign readStage_counterTwoPixelStream_ready = (! readStage_counterTwoPixelStream_rValid);
  assign readStage_counterTwoPixelStream_s2mPipe_valid = (readStage_counterTwoPixelStream_valid || readStage_counterTwoPixelStream_rValid);
  assign readStage_counterTwoPixelStream_s2mPipe_payload = (readStage_counterTwoPixelStream_rValid ? readStage_counterTwoPixelStream_rData : readStage_counterTwoPixelStream_payload);
  always @(*) begin
    readStage_counterTwoPixelStream_s2mPipe_ready = compareStage_counterTwoPixelStream_ready;
    if(when_Stream_l368_31) begin
      readStage_counterTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_31 = (! compareStage_counterTwoPixelStream_valid);
  assign compareStage_counterTwoPixelStream_valid = readStage_counterTwoPixelStream_s2mPipe_rValid;
  assign compareStage_counterTwoPixelStream_payload = readStage_counterTwoPixelStream_s2mPipe_rData;
  assign readStage_mainThreePixelStream_ready = (! readStage_mainThreePixelStream_rValid);
  assign readStage_mainThreePixelStream_s2mPipe_valid = (readStage_mainThreePixelStream_valid || readStage_mainThreePixelStream_rValid);
  assign readStage_mainThreePixelStream_s2mPipe_payload = (readStage_mainThreePixelStream_rValid ? readStage_mainThreePixelStream_rData : readStage_mainThreePixelStream_payload);
  always @(*) begin
    readStage_mainThreePixelStream_s2mPipe_ready = compareStage_mainThreePixelStream_ready;
    if(when_Stream_l368_32) begin
      readStage_mainThreePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_32 = (! compareStage_mainThreePixelStream_valid);
  assign compareStage_mainThreePixelStream_valid = readStage_mainThreePixelStream_s2mPipe_rValid;
  assign compareStage_mainThreePixelStream_payload = readStage_mainThreePixelStream_s2mPipe_rData;
  assign readStage_counterThreePixelStream_ready = (! readStage_counterThreePixelStream_rValid);
  assign readStage_counterThreePixelStream_s2mPipe_valid = (readStage_counterThreePixelStream_valid || readStage_counterThreePixelStream_rValid);
  assign readStage_counterThreePixelStream_s2mPipe_payload = (readStage_counterThreePixelStream_rValid ? readStage_counterThreePixelStream_rData : readStage_counterThreePixelStream_payload);
  always @(*) begin
    readStage_counterThreePixelStream_s2mPipe_ready = compareStage_counterThreePixelStream_ready;
    if(when_Stream_l368_33) begin
      readStage_counterThreePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_33 = (! compareStage_counterThreePixelStream_valid);
  assign compareStage_counterThreePixelStream_valid = readStage_counterThreePixelStream_s2mPipe_rValid;
  assign compareStage_counterThreePixelStream_payload = readStage_counterThreePixelStream_s2mPipe_rData;
  assign readStage_mainOneValidStream_ready = (! readStage_mainOneValidStream_rValid);
  assign readStage_mainOneValidStream_s2mPipe_valid = (readStage_mainOneValidStream_valid || readStage_mainOneValidStream_rValid);
  assign readStage_mainOneValidStream_s2mPipe_payload = (readStage_mainOneValidStream_rValid ? readStage_mainOneValidStream_rData : readStage_mainOneValidStream_payload);
  always @(*) begin
    readStage_mainOneValidStream_s2mPipe_ready = compareStage_mainOneValidStream_ready;
    if(when_Stream_l368_34) begin
      readStage_mainOneValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_34 = (! compareStage_mainOneValidStream_valid);
  assign compareStage_mainOneValidStream_valid = readStage_mainOneValidStream_s2mPipe_rValid;
  assign compareStage_mainOneValidStream_payload = readStage_mainOneValidStream_s2mPipe_rData;
  assign readStage_counterOneValidStream_ready = (! readStage_counterOneValidStream_rValid);
  assign readStage_counterOneValidStream_s2mPipe_valid = (readStage_counterOneValidStream_valid || readStage_counterOneValidStream_rValid);
  assign readStage_counterOneValidStream_s2mPipe_payload = (readStage_counterOneValidStream_rValid ? readStage_counterOneValidStream_rData : readStage_counterOneValidStream_payload);
  always @(*) begin
    readStage_counterOneValidStream_s2mPipe_ready = compareStage_counterOneValidStream_ready;
    if(when_Stream_l368_35) begin
      readStage_counterOneValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_35 = (! compareStage_counterOneValidStream_valid);
  assign compareStage_counterOneValidStream_valid = readStage_counterOneValidStream_s2mPipe_rValid;
  assign compareStage_counterOneValidStream_payload = readStage_counterOneValidStream_s2mPipe_rData;
  assign readStage_mainTwoValidStream_ready = (! readStage_mainTwoValidStream_rValid);
  assign readStage_mainTwoValidStream_s2mPipe_valid = (readStage_mainTwoValidStream_valid || readStage_mainTwoValidStream_rValid);
  assign readStage_mainTwoValidStream_s2mPipe_payload = (readStage_mainTwoValidStream_rValid ? readStage_mainTwoValidStream_rData : readStage_mainTwoValidStream_payload);
  always @(*) begin
    readStage_mainTwoValidStream_s2mPipe_ready = compareStage_mainTwoValidStream_ready;
    if(when_Stream_l368_36) begin
      readStage_mainTwoValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_36 = (! compareStage_mainTwoValidStream_valid);
  assign compareStage_mainTwoValidStream_valid = readStage_mainTwoValidStream_s2mPipe_rValid;
  assign compareStage_mainTwoValidStream_payload = readStage_mainTwoValidStream_s2mPipe_rData;
  assign readStage_counterTwoValidStream_ready = (! readStage_counterTwoValidStream_rValid);
  assign readStage_counterTwoValidStream_s2mPipe_valid = (readStage_counterTwoValidStream_valid || readStage_counterTwoValidStream_rValid);
  assign readStage_counterTwoValidStream_s2mPipe_payload = (readStage_counterTwoValidStream_rValid ? readStage_counterTwoValidStream_rData : readStage_counterTwoValidStream_payload);
  always @(*) begin
    readStage_counterTwoValidStream_s2mPipe_ready = compareStage_counterTwoValidStream_ready;
    if(when_Stream_l368_37) begin
      readStage_counterTwoValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_37 = (! compareStage_counterTwoValidStream_valid);
  assign compareStage_counterTwoValidStream_valid = readStage_counterTwoValidStream_s2mPipe_rValid;
  assign compareStage_counterTwoValidStream_payload = readStage_counterTwoValidStream_s2mPipe_rData;
  assign readStage_mainThreeValidStream_ready = (! readStage_mainThreeValidStream_rValid);
  assign readStage_mainThreeValidStream_s2mPipe_valid = (readStage_mainThreeValidStream_valid || readStage_mainThreeValidStream_rValid);
  assign readStage_mainThreeValidStream_s2mPipe_payload = (readStage_mainThreeValidStream_rValid ? readStage_mainThreeValidStream_rData : readStage_mainThreeValidStream_payload);
  always @(*) begin
    readStage_mainThreeValidStream_s2mPipe_ready = compareStage_mainThreeValidStream_ready;
    if(when_Stream_l368_38) begin
      readStage_mainThreeValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_38 = (! compareStage_mainThreeValidStream_valid);
  assign compareStage_mainThreeValidStream_valid = readStage_mainThreeValidStream_s2mPipe_rValid;
  assign compareStage_mainThreeValidStream_payload = readStage_mainThreeValidStream_s2mPipe_rData;
  assign readStage_counterThreeValidStream_ready = (! readStage_counterThreeValidStream_rValid);
  assign readStage_counterThreeValidStream_s2mPipe_valid = (readStage_counterThreeValidStream_valid || readStage_counterThreeValidStream_rValid);
  assign readStage_counterThreeValidStream_s2mPipe_payload = (readStage_counterThreeValidStream_rValid ? readStage_counterThreeValidStream_rData : readStage_counterThreeValidStream_payload);
  always @(*) begin
    readStage_counterThreeValidStream_s2mPipe_ready = compareStage_counterThreeValidStream_ready;
    if(when_Stream_l368_39) begin
      readStage_counterThreeValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_39 = (! compareStage_counterThreeValidStream_valid);
  assign compareStage_counterThreeValidStream_valid = readStage_counterThreeValidStream_s2mPipe_rValid;
  assign compareStage_counterThreeValidStream_payload = readStage_counterThreeValidStream_s2mPipe_rData;
  always @(*) begin
    CICC1851_readStage_controlPipe_translated_payload_mainCompare = readStage_controlPipe_payload_mainCompare;
    if(!readStage_controlPipe_payload_finalResult) begin
      if(when_SuperResolutionPart3_l415) begin
        if(when_SuperResolutionPart3_l422) begin
          if(readStage_controlPipe_payload_firstRow) begin
            if(when_SuperResolutionPart3_l432) begin
              CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l449) begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l463) begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
              end
            end
          end
        end else begin
          if(readStage_controlPipe_payload_lastRow) begin
            if(when_SuperResolutionPart3_l477) begin
              CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
            end
          end else begin
            if(when_SuperResolutionPart3_l490) begin
              CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
            end
          end
        end
      end else begin
        if(when_SuperResolutionPart3_l496) begin
          if(when_SuperResolutionPart3_l502) begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l511) begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l524) begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
              end
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l539) begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l552) begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
              end
            end
          end
        end else begin
          if(when_SuperResolutionPart3_l564) begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l573) begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l586) begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
              end
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l601) begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l614) begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
              end
            end
          end
        end
      end
    end
  end

  always @(*) begin
    CICC1851_readStage_controlPipe_translated_payload_counterCompare = readStage_controlPipe_payload_counterCompare;
    if(!readStage_controlPipe_payload_finalResult) begin
      if(when_SuperResolutionPart3_l415) begin
        if(when_SuperResolutionPart3_l422) begin
          if(readStage_controlPipe_payload_firstRow) begin
            if(when_SuperResolutionPart3_l432) begin
              CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l449) begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l465) begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
              end
            end
          end
        end else begin
          if(readStage_controlPipe_payload_lastRow) begin
            if(when_SuperResolutionPart3_l477) begin
              CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
            end
          end else begin
            if(when_SuperResolutionPart3_l492) begin
              CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
            end
          end
        end
      end else begin
        if(when_SuperResolutionPart3_l496) begin
          if(when_SuperResolutionPart3_l502) begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l511) begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l526) begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
              end
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l539) begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l554) begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
              end
            end
          end
        end else begin
          if(when_SuperResolutionPart3_l564) begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l573) begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l588) begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
              end
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l601) begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l616) begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
              end
            end
          end
        end
      end
    end
  end

  always @(*) begin
    CICC1851_readStage_controlPipe_translated_payload_horizontalCompare = readStage_controlPipe_payload_horizontalCompare;
    if(!readStage_controlPipe_payload_finalResult) begin
      if(when_SuperResolutionPart3_l415) begin
        if(when_SuperResolutionPart3_l419) begin
          CICC1851_readStage_controlPipe_translated_payload_horizontalCompare = 1'b1;
        end else begin
          CICC1851_readStage_controlPipe_translated_payload_horizontalCompare = 1'b0;
        end
      end else begin
        if(when_SuperResolutionPart3_l496) begin
          if(when_SuperResolutionPart3_l500) begin
            CICC1851_readStage_controlPipe_translated_payload_horizontalCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_horizontalCompare = 1'b0;
          end
        end else begin
          if(when_SuperResolutionPart3_l562) begin
            CICC1851_readStage_controlPipe_translated_payload_horizontalCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_horizontalCompare = 1'b0;
          end
        end
      end
    end
  end

  always @(*) begin
    CICC1851_readStage_controlPipe_translated_payload_verticalCompare = readStage_controlPipe_payload_verticalCompare;
    if(readStage_controlPipe_payload_finalResult) begin
      if(when_SuperResolutionPart3_l342) begin
        CICC1851_readStage_controlPipe_translated_payload_verticalCompare = 1'b1;
      end else begin
        if(when_SuperResolutionPart3_l344) begin
          if(when_SuperResolutionPart3_l345) begin
            CICC1851_readStage_controlPipe_translated_payload_verticalCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_verticalCompare = 1'b0;
          end
        end else begin
          if(when_SuperResolutionPart3_l347) begin
            if(when_SuperResolutionPart3_l348) begin
              CICC1851_readStage_controlPipe_translated_payload_verticalCompare = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_verticalCompare = 1'b0;
            end
          end else begin
            if(when_SuperResolutionPart3_l351) begin
              CICC1851_readStage_controlPipe_translated_payload_verticalCompare = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_verticalCompare = 1'b0;
            end
          end
        end
      end
    end
  end

  always @(*) begin
    CICC1851_readStage_controlPipe_translated_payload_horizontalDirectionValid = readStage_controlPipe_payload_horizontalDirectionValid;
    if(!readStage_controlPipe_payload_finalResult) begin
      if(when_SuperResolutionPart3_l415) begin
        if(when_SuperResolutionPart3_l416) begin
          CICC1851_readStage_controlPipe_translated_payload_horizontalDirectionValid = 1'b1;
        end else begin
          CICC1851_readStage_controlPipe_translated_payload_horizontalDirectionValid = 1'b0;
        end
      end else begin
        if(when_SuperResolutionPart3_l496) begin
          if(when_SuperResolutionPart3_l497) begin
            CICC1851_readStage_controlPipe_translated_payload_horizontalDirectionValid = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_horizontalDirectionValid = 1'b0;
          end
        end else begin
          if(when_SuperResolutionPart3_l559) begin
            CICC1851_readStage_controlPipe_translated_payload_horizontalDirectionValid = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_horizontalDirectionValid = 1'b0;
          end
        end
      end
    end
  end

  always @(*) begin
    CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = readStage_controlPipe_payload_verticalDirectionValid;
    if(readStage_controlPipe_payload_finalResult) begin
      if(when_SuperResolutionPart3_l356) begin
        if(when_SuperResolutionPart3_l357) begin
          if(readStage_controlPipe_payload_firstRow) begin
            if(readStage_mainTwoValidStream_payload) begin
              CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b0;
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(readStage_mainThreeValidStream_payload) begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l365) begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b0;
              end
            end
          end
        end else begin
          if(readStage_controlPipe_payload_lastRow) begin
            if(readStage_mainTwoValidStream_payload) begin
              CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b0;
            end
          end else begin
            if(when_SuperResolutionPart3_l373) begin
              CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b0;
            end
          end
        end
      end else begin
        if(when_SuperResolutionPart3_l377) begin
          if(when_SuperResolutionPart3_l378) begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(readStage_mainThreeValidStream_payload) begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l383) begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b0;
              end
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(readStage_mainOneValidStream_payload) begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l391) begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b0;
              end
            end
          end
        end else begin
          if(when_SuperResolutionPart3_l396) begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(readStage_mainTwoValidStream_payload) begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l401) begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b0;
              end
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(readStage_mainOneValidStream_payload) begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l409) begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid = 1'b0;
              end
            end
          end
        end
      end
    end
  end

  always @(*) begin
    CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = readStage_controlPipe_payload_mainDirectionValid;
    if(!readStage_controlPipe_payload_finalResult) begin
      if(when_SuperResolutionPart3_l415) begin
        if(when_SuperResolutionPart3_l422) begin
          if(readStage_controlPipe_payload_firstRow) begin
            if(when_SuperResolutionPart3_l424) begin
              CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b0;
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l441) begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l458) begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b0;
              end
            end
          end
        end else begin
          if(readStage_controlPipe_payload_lastRow) begin
            if(when_SuperResolutionPart3_l470) begin
              CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b0;
            end
          end else begin
            if(when_SuperResolutionPart3_l485) begin
              CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b0;
            end
          end
        end
      end else begin
        if(when_SuperResolutionPart3_l496) begin
          if(when_SuperResolutionPart3_l502) begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l504) begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l519) begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b0;
              end
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l531) begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l547) begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b0;
              end
            end
          end
        end else begin
          if(when_SuperResolutionPart3_l564) begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l566) begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l581) begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b0;
              end
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l593) begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l609) begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid = 1'b0;
              end
            end
          end
        end
      end
    end
  end

  always @(*) begin
    CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = readStage_controlPipe_payload_counterDirectionValid;
    if(!readStage_controlPipe_payload_finalResult) begin
      if(when_SuperResolutionPart3_l415) begin
        if(when_SuperResolutionPart3_l422) begin
          if(readStage_controlPipe_payload_firstRow) begin
            if(when_SuperResolutionPart3_l424) begin
              CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b0;
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l441) begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l460) begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b0;
              end
            end
          end
        end else begin
          if(readStage_controlPipe_payload_lastRow) begin
            if(when_SuperResolutionPart3_l470) begin
              CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b0;
            end
          end else begin
            if(when_SuperResolutionPart3_l487) begin
              CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b1;
            end else begin
              CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b0;
            end
          end
        end
      end else begin
        if(when_SuperResolutionPart3_l496) begin
          if(when_SuperResolutionPart3_l502) begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l504) begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l521) begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b0;
              end
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l531) begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l549) begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b0;
              end
            end
          end
        end else begin
          if(when_SuperResolutionPart3_l564) begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l566) begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l583) begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b0;
              end
            end
          end else begin
            if(readStage_controlPipe_payload_lastRow) begin
              if(when_SuperResolutionPart3_l593) begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l611) begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b1;
              end else begin
                CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid = 1'b0;
              end
            end
          end
        end
      end
    end
  end

  assign when_SuperResolutionPart3_l342 = (readStage_controlPipe_payload_firstRow || readStage_controlPipe_payload_lastRow);
  assign when_SuperResolutionPart3_l344 = (readStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l345 = (readStage_mainThreePixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart3_l348 = (readStage_mainThreePixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart3_l351 = (readStage_mainTwoPixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart3_l347 = (readStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l356 = (readStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l357 = (readStage_controlPipe_payload_nextPosition == 2'b01);
  assign when_SuperResolutionPart3_l365 = (readStage_mainTwoValidStream_payload && readStage_mainThreeValidStream_payload);
  assign when_SuperResolutionPart3_l373 = (readStage_mainTwoValidStream_payload && readStage_mainThreeValidStream_payload);
  assign when_SuperResolutionPart3_l378 = (readStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l383 = (readStage_mainOneValidStream_payload && readStage_mainThreeValidStream_payload);
  assign when_SuperResolutionPart3_l391 = (readStage_mainOneValidStream_payload && readStage_mainThreeValidStream_payload);
  assign when_SuperResolutionPart3_l396 = (readStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l401 = (readStage_mainOneValidStream_payload && readStage_mainTwoValidStream_payload);
  assign when_SuperResolutionPart3_l409 = (readStage_mainOneValidStream_payload && readStage_mainTwoValidStream_payload);
  assign when_SuperResolutionPart3_l377 = (readStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l415 = (readStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l416 = (readStage_mainOneValidStream_payload && readStage_counterOneValidStream_payload);
  assign when_SuperResolutionPart3_l419 = (readStage_counterOnePixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart3_l422 = (readStage_controlPipe_payload_nextPosition == 2'b01);
  assign when_SuperResolutionPart3_l424 = (readStage_mainTwoValidStream_payload && readStage_counterTwoValidStream_payload);
  assign when_SuperResolutionPart3_l432 = (readStage_counterTwoPixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart3_l441 = (readStage_mainThreeValidStream_payload && readStage_counterThreeValidStream_payload);
  assign when_SuperResolutionPart3_l449 = (readStage_counterThreePixelStream_payload <= readStage_mainThreePixelStream_payload);
  assign when_SuperResolutionPart3_l458 = (readStage_mainThreeValidStream_payload && readStage_counterTwoValidStream_payload);
  assign when_SuperResolutionPart3_l460 = (readStage_mainTwoValidStream_payload && readStage_counterThreeValidStream_payload);
  assign when_SuperResolutionPart3_l463 = (readStage_counterTwoPixelStream_payload <= readStage_mainThreePixelStream_payload);
  assign when_SuperResolutionPart3_l465 = (readStage_counterThreePixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart3_l470 = (readStage_mainTwoValidStream_payload && readStage_counterTwoValidStream_payload);
  assign when_SuperResolutionPart3_l477 = (readStage_counterTwoPixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart3_l485 = (readStage_mainTwoValidStream_payload && readStage_counterThreeValidStream_payload);
  assign when_SuperResolutionPart3_l487 = (readStage_mainThreeValidStream_payload && readStage_counterTwoValidStream_payload);
  assign when_SuperResolutionPart3_l490 = (readStage_counterThreePixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart3_l492 = (readStage_counterTwoPixelStream_payload <= readStage_mainThreePixelStream_payload);
  assign when_SuperResolutionPart3_l497 = (readStage_mainTwoValidStream_payload && readStage_counterTwoValidStream_payload);
  assign when_SuperResolutionPart3_l500 = (readStage_counterTwoPixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart3_l502 = (readStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l504 = (readStage_mainThreeValidStream_payload && readStage_counterThreeValidStream_payload);
  assign when_SuperResolutionPart3_l511 = (readStage_counterThreePixelStream_payload <= readStage_mainThreePixelStream_payload);
  assign when_SuperResolutionPart3_l519 = (readStage_mainThreeValidStream_payload && readStage_counterOneValidStream_payload);
  assign when_SuperResolutionPart3_l521 = (readStage_mainOneValidStream_payload && readStage_counterThreeValidStream_payload);
  assign when_SuperResolutionPart3_l524 = (readStage_counterOnePixelStream_payload <= readStage_mainThreePixelStream_payload);
  assign when_SuperResolutionPart3_l526 = (readStage_counterThreePixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart3_l531 = (readStage_mainOneValidStream_payload && readStage_counterOneValidStream_payload);
  assign when_SuperResolutionPart3_l539 = (readStage_counterOnePixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart3_l547 = (readStage_mainOneValidStream_payload && readStage_counterThreeValidStream_payload);
  assign when_SuperResolutionPart3_l549 = (readStage_mainThreeValidStream_payload && readStage_counterOneValidStream_payload);
  assign when_SuperResolutionPart3_l552 = (readStage_counterThreePixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart3_l554 = (readStage_counterOnePixelStream_payload <= readStage_mainThreePixelStream_payload);
  assign when_SuperResolutionPart3_l559 = (readStage_mainThreeValidStream_payload && readStage_counterThreeValidStream_payload);
  assign when_SuperResolutionPart3_l562 = (readStage_counterThreePixelStream_payload <= readStage_mainThreePixelStream_payload);
  assign when_SuperResolutionPart3_l564 = (readStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l566 = (readStage_mainTwoValidStream_payload && readStage_counterTwoValidStream_payload);
  assign when_SuperResolutionPart3_l573 = (readStage_counterTwoPixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart3_l581 = (readStage_mainTwoValidStream_payload && readStage_counterOneValidStream_payload);
  assign when_SuperResolutionPart3_l583 = (readStage_mainOneValidStream_payload && readStage_counterTwoValidStream_payload);
  assign when_SuperResolutionPart3_l586 = (readStage_counterOnePixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart3_l588 = (readStage_counterTwoPixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart3_l593 = (readStage_mainOneValidStream_payload && readStage_counterOneValidStream_payload);
  assign when_SuperResolutionPart3_l601 = (readStage_counterOnePixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart3_l609 = (readStage_mainOneValidStream_payload && readStage_counterTwoValidStream_payload);
  assign when_SuperResolutionPart3_l611 = (readStage_mainTwoValidStream_payload && readStage_counterOneValidStream_payload);
  assign when_SuperResolutionPart3_l614 = (readStage_counterTwoPixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart3_l616 = (readStage_counterOnePixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart3_l496 = (readStage_controlPipe_payload_currentPosition == 2'b01);
  assign readStage_controlPipe_translated_valid = readStage_controlPipe_valid;
  assign readStage_controlPipe_ready = readStage_controlPipe_translated_ready;
  assign readStage_controlPipe_translated_payload_frameStart = readStage_controlPipe_payload_frameStart;
  assign readStage_controlPipe_translated_payload_rowEnd = readStage_controlPipe_payload_rowEnd;
  assign readStage_controlPipe_translated_payload_pipeValid = readStage_controlPipe_payload_pipeValid;
  assign readStage_controlPipe_translated_payload_firstRow = readStage_controlPipe_payload_firstRow;
  assign readStage_controlPipe_translated_payload_lastRow = readStage_controlPipe_payload_lastRow;
  assign readStage_controlPipe_translated_payload_finalResult = readStage_controlPipe_payload_finalResult;
  assign readStage_controlPipe_translated_payload_mainCompare = CICC1851_readStage_controlPipe_translated_payload_mainCompare;
  assign readStage_controlPipe_translated_payload_counterCompare = CICC1851_readStage_controlPipe_translated_payload_counterCompare;
  assign readStage_controlPipe_translated_payload_horizontalCompare = CICC1851_readStage_controlPipe_translated_payload_horizontalCompare;
  assign readStage_controlPipe_translated_payload_verticalCompare = CICC1851_readStage_controlPipe_translated_payload_verticalCompare;
  assign readStage_controlPipe_translated_payload_mainDiff = readStage_controlPipe_payload_mainDiff;
  assign readStage_controlPipe_translated_payload_counterDiff = readStage_controlPipe_payload_counterDiff;
  assign readStage_controlPipe_translated_payload_horizontalDiff = readStage_controlPipe_payload_horizontalDiff;
  assign readStage_controlPipe_translated_payload_verticalDiff = readStage_controlPipe_payload_verticalDiff;
  assign readStage_controlPipe_translated_payload_isHorizontalMin = readStage_controlPipe_payload_isHorizontalMin;
  assign readStage_controlPipe_translated_payload_minDiff = readStage_controlPipe_payload_minDiff;
  assign readStage_controlPipe_translated_payload_currentPosition = readStage_controlPipe_payload_currentPosition;
  assign readStage_controlPipe_translated_payload_nextPosition = readStage_controlPipe_payload_nextPosition;
  assign readStage_controlPipe_translated_payload_horizontalDirectionValid = CICC1851_readStage_controlPipe_translated_payload_horizontalDirectionValid;
  assign readStage_controlPipe_translated_payload_verticalDirectionValid = CICC1851_readStage_controlPipe_translated_payload_verticalDirectionValid;
  assign readStage_controlPipe_translated_payload_mainDirectionValid = CICC1851_readStage_controlPipe_translated_payload_mainDirectionValid;
  assign readStage_controlPipe_translated_payload_counterDirectionValid = CICC1851_readStage_controlPipe_translated_payload_counterDirectionValid;
  assign readStage_controlPipe_translated_payload_inValidMinDiff = readStage_controlPipe_payload_inValidMinDiff;
  assign readStage_controlPipe_translated_ready = (! readStage_controlPipe_translated_rValid);
  assign readStage_controlPipe_translated_s2mPipe_valid = (readStage_controlPipe_translated_valid || readStage_controlPipe_translated_rValid);
  assign readStage_controlPipe_translated_s2mPipe_payload_frameStart = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_frameStart : readStage_controlPipe_translated_payload_frameStart);
  assign readStage_controlPipe_translated_s2mPipe_payload_rowEnd = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_rowEnd : readStage_controlPipe_translated_payload_rowEnd);
  assign readStage_controlPipe_translated_s2mPipe_payload_pipeValid = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_pipeValid : readStage_controlPipe_translated_payload_pipeValid);
  assign readStage_controlPipe_translated_s2mPipe_payload_firstRow = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_firstRow : readStage_controlPipe_translated_payload_firstRow);
  assign readStage_controlPipe_translated_s2mPipe_payload_lastRow = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_lastRow : readStage_controlPipe_translated_payload_lastRow);
  assign readStage_controlPipe_translated_s2mPipe_payload_finalResult = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_finalResult : readStage_controlPipe_translated_payload_finalResult);
  assign readStage_controlPipe_translated_s2mPipe_payload_mainCompare = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_mainCompare : readStage_controlPipe_translated_payload_mainCompare);
  assign readStage_controlPipe_translated_s2mPipe_payload_counterCompare = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_counterCompare : readStage_controlPipe_translated_payload_counterCompare);
  assign readStage_controlPipe_translated_s2mPipe_payload_horizontalCompare = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_horizontalCompare : readStage_controlPipe_translated_payload_horizontalCompare);
  assign readStage_controlPipe_translated_s2mPipe_payload_verticalCompare = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_verticalCompare : readStage_controlPipe_translated_payload_verticalCompare);
  assign readStage_controlPipe_translated_s2mPipe_payload_mainDiff = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_mainDiff : readStage_controlPipe_translated_payload_mainDiff);
  assign readStage_controlPipe_translated_s2mPipe_payload_counterDiff = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_counterDiff : readStage_controlPipe_translated_payload_counterDiff);
  assign readStage_controlPipe_translated_s2mPipe_payload_horizontalDiff = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_horizontalDiff : readStage_controlPipe_translated_payload_horizontalDiff);
  assign readStage_controlPipe_translated_s2mPipe_payload_verticalDiff = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_verticalDiff : readStage_controlPipe_translated_payload_verticalDiff);
  assign readStage_controlPipe_translated_s2mPipe_payload_isHorizontalMin = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_isHorizontalMin : readStage_controlPipe_translated_payload_isHorizontalMin);
  assign readStage_controlPipe_translated_s2mPipe_payload_minDiff = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_minDiff : readStage_controlPipe_translated_payload_minDiff);
  assign readStage_controlPipe_translated_s2mPipe_payload_currentPosition = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_currentPosition : readStage_controlPipe_translated_payload_currentPosition);
  assign readStage_controlPipe_translated_s2mPipe_payload_nextPosition = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_nextPosition : readStage_controlPipe_translated_payload_nextPosition);
  assign readStage_controlPipe_translated_s2mPipe_payload_horizontalDirectionValid = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_horizontalDirectionValid : readStage_controlPipe_translated_payload_horizontalDirectionValid);
  assign readStage_controlPipe_translated_s2mPipe_payload_verticalDirectionValid = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_verticalDirectionValid : readStage_controlPipe_translated_payload_verticalDirectionValid);
  assign readStage_controlPipe_translated_s2mPipe_payload_mainDirectionValid = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_mainDirectionValid : readStage_controlPipe_translated_payload_mainDirectionValid);
  assign readStage_controlPipe_translated_s2mPipe_payload_counterDirectionValid = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_counterDirectionValid : readStage_controlPipe_translated_payload_counterDirectionValid);
  assign readStage_controlPipe_translated_s2mPipe_payload_inValidMinDiff = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_inValidMinDiff : readStage_controlPipe_translated_payload_inValidMinDiff);
  always @(*) begin
    readStage_controlPipe_translated_s2mPipe_ready = compareStage_controlPipe_ready;
    if(when_Stream_l368_40) begin
      readStage_controlPipe_translated_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_40 = (! compareStage_controlPipe_valid);
  assign compareStage_controlPipe_valid = readStage_controlPipe_translated_s2mPipe_rValid;
  assign compareStage_controlPipe_payload_frameStart = readStage_controlPipe_translated_s2mPipe_rData_frameStart;
  assign compareStage_controlPipe_payload_rowEnd = readStage_controlPipe_translated_s2mPipe_rData_rowEnd;
  assign compareStage_controlPipe_payload_pipeValid = readStage_controlPipe_translated_s2mPipe_rData_pipeValid;
  assign compareStage_controlPipe_payload_firstRow = readStage_controlPipe_translated_s2mPipe_rData_firstRow;
  assign compareStage_controlPipe_payload_lastRow = readStage_controlPipe_translated_s2mPipe_rData_lastRow;
  assign compareStage_controlPipe_payload_finalResult = readStage_controlPipe_translated_s2mPipe_rData_finalResult;
  assign compareStage_controlPipe_payload_mainCompare = readStage_controlPipe_translated_s2mPipe_rData_mainCompare;
  assign compareStage_controlPipe_payload_counterCompare = readStage_controlPipe_translated_s2mPipe_rData_counterCompare;
  assign compareStage_controlPipe_payload_horizontalCompare = readStage_controlPipe_translated_s2mPipe_rData_horizontalCompare;
  assign compareStage_controlPipe_payload_verticalCompare = readStage_controlPipe_translated_s2mPipe_rData_verticalCompare;
  assign compareStage_controlPipe_payload_mainDiff = readStage_controlPipe_translated_s2mPipe_rData_mainDiff;
  assign compareStage_controlPipe_payload_counterDiff = readStage_controlPipe_translated_s2mPipe_rData_counterDiff;
  assign compareStage_controlPipe_payload_horizontalDiff = readStage_controlPipe_translated_s2mPipe_rData_horizontalDiff;
  assign compareStage_controlPipe_payload_verticalDiff = readStage_controlPipe_translated_s2mPipe_rData_verticalDiff;
  assign compareStage_controlPipe_payload_isHorizontalMin = readStage_controlPipe_translated_s2mPipe_rData_isHorizontalMin;
  assign compareStage_controlPipe_payload_minDiff = readStage_controlPipe_translated_s2mPipe_rData_minDiff;
  assign compareStage_controlPipe_payload_currentPosition = readStage_controlPipe_translated_s2mPipe_rData_currentPosition;
  assign compareStage_controlPipe_payload_nextPosition = readStage_controlPipe_translated_s2mPipe_rData_nextPosition;
  assign compareStage_controlPipe_payload_horizontalDirectionValid = readStage_controlPipe_translated_s2mPipe_rData_horizontalDirectionValid;
  assign compareStage_controlPipe_payload_verticalDirectionValid = readStage_controlPipe_translated_s2mPipe_rData_verticalDirectionValid;
  assign compareStage_controlPipe_payload_mainDirectionValid = readStage_controlPipe_translated_s2mPipe_rData_mainDirectionValid;
  assign compareStage_controlPipe_payload_counterDirectionValid = readStage_controlPipe_translated_s2mPipe_rData_counterDirectionValid;
  assign compareStage_controlPipe_payload_inValidMinDiff = readStage_controlPipe_translated_s2mPipe_rData_inValidMinDiff;
  assign compareStage_mainOnePixelStream_ready = (! compareStage_mainOnePixelStream_rValid);
  assign compareStage_mainOnePixelStream_s2mPipe_valid = (compareStage_mainOnePixelStream_valid || compareStage_mainOnePixelStream_rValid);
  assign compareStage_mainOnePixelStream_s2mPipe_payload = (compareStage_mainOnePixelStream_rValid ? compareStage_mainOnePixelStream_rData : compareStage_mainOnePixelStream_payload);
  always @(*) begin
    compareStage_mainOnePixelStream_s2mPipe_ready = diffStage_mainOnePixelStream_ready;
    if(when_Stream_l368_41) begin
      compareStage_mainOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_41 = (! diffStage_mainOnePixelStream_valid);
  assign diffStage_mainOnePixelStream_valid = compareStage_mainOnePixelStream_s2mPipe_rValid;
  assign diffStage_mainOnePixelStream_payload = compareStage_mainOnePixelStream_s2mPipe_rData;
  assign compareStage_counterOnePixelStream_ready = (! compareStage_counterOnePixelStream_rValid);
  assign compareStage_counterOnePixelStream_s2mPipe_valid = (compareStage_counterOnePixelStream_valid || compareStage_counterOnePixelStream_rValid);
  assign compareStage_counterOnePixelStream_s2mPipe_payload = (compareStage_counterOnePixelStream_rValid ? compareStage_counterOnePixelStream_rData : compareStage_counterOnePixelStream_payload);
  always @(*) begin
    compareStage_counterOnePixelStream_s2mPipe_ready = diffStage_counterOnePixelStream_ready;
    if(when_Stream_l368_42) begin
      compareStage_counterOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_42 = (! diffStage_counterOnePixelStream_valid);
  assign diffStage_counterOnePixelStream_valid = compareStage_counterOnePixelStream_s2mPipe_rValid;
  assign diffStage_counterOnePixelStream_payload = compareStage_counterOnePixelStream_s2mPipe_rData;
  assign compareStage_mainTwoPixelStream_ready = (! compareStage_mainTwoPixelStream_rValid);
  assign compareStage_mainTwoPixelStream_s2mPipe_valid = (compareStage_mainTwoPixelStream_valid || compareStage_mainTwoPixelStream_rValid);
  assign compareStage_mainTwoPixelStream_s2mPipe_payload = (compareStage_mainTwoPixelStream_rValid ? compareStage_mainTwoPixelStream_rData : compareStage_mainTwoPixelStream_payload);
  always @(*) begin
    compareStage_mainTwoPixelStream_s2mPipe_ready = diffStage_mainTwoPixelStream_ready;
    if(when_Stream_l368_43) begin
      compareStage_mainTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_43 = (! diffStage_mainTwoPixelStream_valid);
  assign diffStage_mainTwoPixelStream_valid = compareStage_mainTwoPixelStream_s2mPipe_rValid;
  assign diffStage_mainTwoPixelStream_payload = compareStage_mainTwoPixelStream_s2mPipe_rData;
  assign compareStage_counterTwoPixelStream_ready = (! compareStage_counterTwoPixelStream_rValid);
  assign compareStage_counterTwoPixelStream_s2mPipe_valid = (compareStage_counterTwoPixelStream_valid || compareStage_counterTwoPixelStream_rValid);
  assign compareStage_counterTwoPixelStream_s2mPipe_payload = (compareStage_counterTwoPixelStream_rValid ? compareStage_counterTwoPixelStream_rData : compareStage_counterTwoPixelStream_payload);
  always @(*) begin
    compareStage_counterTwoPixelStream_s2mPipe_ready = diffStage_counterTwoPixelStream_ready;
    if(when_Stream_l368_44) begin
      compareStage_counterTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_44 = (! diffStage_counterTwoPixelStream_valid);
  assign diffStage_counterTwoPixelStream_valid = compareStage_counterTwoPixelStream_s2mPipe_rValid;
  assign diffStage_counterTwoPixelStream_payload = compareStage_counterTwoPixelStream_s2mPipe_rData;
  assign compareStage_mainThreePixelStream_ready = (! compareStage_mainThreePixelStream_rValid);
  assign compareStage_mainThreePixelStream_s2mPipe_valid = (compareStage_mainThreePixelStream_valid || compareStage_mainThreePixelStream_rValid);
  assign compareStage_mainThreePixelStream_s2mPipe_payload = (compareStage_mainThreePixelStream_rValid ? compareStage_mainThreePixelStream_rData : compareStage_mainThreePixelStream_payload);
  always @(*) begin
    compareStage_mainThreePixelStream_s2mPipe_ready = diffStage_mainThreePixelStream_ready;
    if(when_Stream_l368_45) begin
      compareStage_mainThreePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_45 = (! diffStage_mainThreePixelStream_valid);
  assign diffStage_mainThreePixelStream_valid = compareStage_mainThreePixelStream_s2mPipe_rValid;
  assign diffStage_mainThreePixelStream_payload = compareStage_mainThreePixelStream_s2mPipe_rData;
  assign compareStage_counterThreePixelStream_ready = (! compareStage_counterThreePixelStream_rValid);
  assign compareStage_counterThreePixelStream_s2mPipe_valid = (compareStage_counterThreePixelStream_valid || compareStage_counterThreePixelStream_rValid);
  assign compareStage_counterThreePixelStream_s2mPipe_payload = (compareStage_counterThreePixelStream_rValid ? compareStage_counterThreePixelStream_rData : compareStage_counterThreePixelStream_payload);
  always @(*) begin
    compareStage_counterThreePixelStream_s2mPipe_ready = diffStage_counterThreePixelStream_ready;
    if(when_Stream_l368_46) begin
      compareStage_counterThreePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_46 = (! diffStage_counterThreePixelStream_valid);
  assign diffStage_counterThreePixelStream_valid = compareStage_counterThreePixelStream_s2mPipe_rValid;
  assign diffStage_counterThreePixelStream_payload = compareStage_counterThreePixelStream_s2mPipe_rData;
  assign compareStage_mainOneValidStream_ready = (! compareStage_mainOneValidStream_rValid);
  assign compareStage_mainOneValidStream_s2mPipe_valid = (compareStage_mainOneValidStream_valid || compareStage_mainOneValidStream_rValid);
  assign compareStage_mainOneValidStream_s2mPipe_payload = (compareStage_mainOneValidStream_rValid ? compareStage_mainOneValidStream_rData : compareStage_mainOneValidStream_payload);
  always @(*) begin
    compareStage_mainOneValidStream_s2mPipe_ready = diffStage_mainOneValidStream_ready;
    if(when_Stream_l368_47) begin
      compareStage_mainOneValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_47 = (! diffStage_mainOneValidStream_valid);
  assign diffStage_mainOneValidStream_valid = compareStage_mainOneValidStream_s2mPipe_rValid;
  assign diffStage_mainOneValidStream_payload = compareStage_mainOneValidStream_s2mPipe_rData;
  assign compareStage_counterOneValidStream_ready = (! compareStage_counterOneValidStream_rValid);
  assign compareStage_counterOneValidStream_s2mPipe_valid = (compareStage_counterOneValidStream_valid || compareStage_counterOneValidStream_rValid);
  assign compareStage_counterOneValidStream_s2mPipe_payload = (compareStage_counterOneValidStream_rValid ? compareStage_counterOneValidStream_rData : compareStage_counterOneValidStream_payload);
  always @(*) begin
    compareStage_counterOneValidStream_s2mPipe_ready = diffStage_counterOneValidStream_ready;
    if(when_Stream_l368_48) begin
      compareStage_counterOneValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_48 = (! diffStage_counterOneValidStream_valid);
  assign diffStage_counterOneValidStream_valid = compareStage_counterOneValidStream_s2mPipe_rValid;
  assign diffStage_counterOneValidStream_payload = compareStage_counterOneValidStream_s2mPipe_rData;
  assign compareStage_mainTwoValidStream_ready = (! compareStage_mainTwoValidStream_rValid);
  assign compareStage_mainTwoValidStream_s2mPipe_valid = (compareStage_mainTwoValidStream_valid || compareStage_mainTwoValidStream_rValid);
  assign compareStage_mainTwoValidStream_s2mPipe_payload = (compareStage_mainTwoValidStream_rValid ? compareStage_mainTwoValidStream_rData : compareStage_mainTwoValidStream_payload);
  always @(*) begin
    compareStage_mainTwoValidStream_s2mPipe_ready = diffStage_mainTwoValidStream_ready;
    if(when_Stream_l368_49) begin
      compareStage_mainTwoValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_49 = (! diffStage_mainTwoValidStream_valid);
  assign diffStage_mainTwoValidStream_valid = compareStage_mainTwoValidStream_s2mPipe_rValid;
  assign diffStage_mainTwoValidStream_payload = compareStage_mainTwoValidStream_s2mPipe_rData;
  assign compareStage_counterTwoValidStream_ready = (! compareStage_counterTwoValidStream_rValid);
  assign compareStage_counterTwoValidStream_s2mPipe_valid = (compareStage_counterTwoValidStream_valid || compareStage_counterTwoValidStream_rValid);
  assign compareStage_counterTwoValidStream_s2mPipe_payload = (compareStage_counterTwoValidStream_rValid ? compareStage_counterTwoValidStream_rData : compareStage_counterTwoValidStream_payload);
  always @(*) begin
    compareStage_counterTwoValidStream_s2mPipe_ready = diffStage_counterTwoValidStream_ready;
    if(when_Stream_l368_50) begin
      compareStage_counterTwoValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_50 = (! diffStage_counterTwoValidStream_valid);
  assign diffStage_counterTwoValidStream_valid = compareStage_counterTwoValidStream_s2mPipe_rValid;
  assign diffStage_counterTwoValidStream_payload = compareStage_counterTwoValidStream_s2mPipe_rData;
  assign compareStage_mainThreeValidStream_ready = (! compareStage_mainThreeValidStream_rValid);
  assign compareStage_mainThreeValidStream_s2mPipe_valid = (compareStage_mainThreeValidStream_valid || compareStage_mainThreeValidStream_rValid);
  assign compareStage_mainThreeValidStream_s2mPipe_payload = (compareStage_mainThreeValidStream_rValid ? compareStage_mainThreeValidStream_rData : compareStage_mainThreeValidStream_payload);
  always @(*) begin
    compareStage_mainThreeValidStream_s2mPipe_ready = diffStage_mainThreeValidStream_ready;
    if(when_Stream_l368_51) begin
      compareStage_mainThreeValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_51 = (! diffStage_mainThreeValidStream_valid);
  assign diffStage_mainThreeValidStream_valid = compareStage_mainThreeValidStream_s2mPipe_rValid;
  assign diffStage_mainThreeValidStream_payload = compareStage_mainThreeValidStream_s2mPipe_rData;
  assign compareStage_counterThreeValidStream_ready = (! compareStage_counterThreeValidStream_rValid);
  assign compareStage_counterThreeValidStream_s2mPipe_valid = (compareStage_counterThreeValidStream_valid || compareStage_counterThreeValidStream_rValid);
  assign compareStage_counterThreeValidStream_s2mPipe_payload = (compareStage_counterThreeValidStream_rValid ? compareStage_counterThreeValidStream_rData : compareStage_counterThreeValidStream_payload);
  always @(*) begin
    compareStage_counterThreeValidStream_s2mPipe_ready = diffStage_counterThreeValidStream_ready;
    if(when_Stream_l368_52) begin
      compareStage_counterThreeValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_52 = (! diffStage_counterThreeValidStream_valid);
  assign diffStage_counterThreeValidStream_valid = compareStage_counterThreeValidStream_s2mPipe_rValid;
  assign diffStage_counterThreeValidStream_payload = compareStage_counterThreeValidStream_s2mPipe_rData;
  always @(*) begin
    CICC1851_compareStage_controlPipe_translated_payload_mainDiff = compareStage_controlPipe_payload_mainDiff;
    if(!compareStage_controlPipe_payload_finalResult) begin
      if(when_SuperResolutionPart3_l661) begin
        if(when_SuperResolutionPart3_l664) begin
          if(compareStage_controlPipe_payload_firstRow) begin
            if(compareStage_controlPipe_payload_mainCompare) begin
              CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterTwoPixelStream_payload);
            end else begin
              CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainTwoPixelStream_payload);
            end
          end else begin
            if(compareStage_controlPipe_payload_lastRow) begin
              if(compareStage_controlPipe_payload_mainCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainThreePixelStream_payload - compareStage_counterThreePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterThreePixelStream_payload - compareStage_mainThreePixelStream_payload);
              end
            end else begin
              if(compareStage_controlPipe_payload_mainCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainThreePixelStream_payload - compareStage_counterTwoPixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainThreePixelStream_payload);
              end
            end
          end
        end else begin
          if(compareStage_controlPipe_payload_lastRow) begin
            if(compareStage_controlPipe_payload_mainCompare) begin
              CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterTwoPixelStream_payload);
            end else begin
              CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainTwoPixelStream_payload);
            end
          end else begin
            if(compareStage_controlPipe_payload_mainCompare) begin
              CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterThreePixelStream_payload);
            end else begin
              CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterThreePixelStream_payload - compareStage_mainTwoPixelStream_payload);
            end
          end
        end
      end else begin
        if(when_SuperResolutionPart3_l694) begin
          if(when_SuperResolutionPart3_l697) begin
            if(compareStage_controlPipe_payload_lastRow) begin
              if(compareStage_controlPipe_payload_mainCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainThreePixelStream_payload - compareStage_counterThreePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterThreePixelStream_payload - compareStage_mainThreePixelStream_payload);
              end
            end else begin
              if(compareStage_controlPipe_payload_mainCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainThreePixelStream_payload - compareStage_counterOnePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterOnePixelStream_payload - compareStage_mainThreePixelStream_payload);
              end
            end
          end else begin
            if(compareStage_controlPipe_payload_lastRow) begin
              if(compareStage_controlPipe_payload_mainCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_counterOnePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterOnePixelStream_payload - compareStage_mainOnePixelStream_payload);
              end
            end else begin
              if(compareStage_controlPipe_payload_mainCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_counterThreePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterThreePixelStream_payload - compareStage_mainOnePixelStream_payload);
              end
            end
          end
        end else begin
          if(when_SuperResolutionPart3_l725) begin
            if(compareStage_controlPipe_payload_lastRow) begin
              if(compareStage_controlPipe_payload_mainCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterTwoPixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainTwoPixelStream_payload);
              end
            end else begin
              if(compareStage_controlPipe_payload_mainCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterOnePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterOnePixelStream_payload - compareStage_mainTwoPixelStream_payload);
              end
            end
          end else begin
            if(compareStage_controlPipe_payload_lastRow) begin
              if(compareStage_controlPipe_payload_mainCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_counterOnePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterOnePixelStream_payload - compareStage_mainOnePixelStream_payload);
              end
            end else begin
              if(compareStage_controlPipe_payload_mainCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_counterTwoPixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainOnePixelStream_payload);
              end
            end
          end
        end
      end
    end
  end

  always @(*) begin
    CICC1851_compareStage_controlPipe_translated_payload_counterDiff = compareStage_controlPipe_payload_counterDiff;
    if(!compareStage_controlPipe_payload_finalResult) begin
      if(when_SuperResolutionPart3_l661) begin
        if(when_SuperResolutionPart3_l664) begin
          if(compareStage_controlPipe_payload_firstRow) begin
            if(compareStage_controlPipe_payload_counterCompare) begin
              CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterTwoPixelStream_payload);
            end else begin
              CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainTwoPixelStream_payload);
            end
          end else begin
            if(compareStage_controlPipe_payload_lastRow) begin
              if(compareStage_controlPipe_payload_counterCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_mainThreePixelStream_payload - compareStage_counterThreePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterThreePixelStream_payload - compareStage_mainThreePixelStream_payload);
              end
            end else begin
              if(compareStage_controlPipe_payload_counterCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterThreePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterThreePixelStream_payload - compareStage_mainTwoPixelStream_payload);
              end
            end
          end
        end else begin
          if(compareStage_controlPipe_payload_lastRow) begin
            if(compareStage_controlPipe_payload_counterCompare) begin
              CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterTwoPixelStream_payload);
            end else begin
              CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainTwoPixelStream_payload);
            end
          end else begin
            if(compareStage_controlPipe_payload_counterCompare) begin
              CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_mainThreePixelStream_payload - compareStage_counterTwoPixelStream_payload);
            end else begin
              CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainThreePixelStream_payload);
            end
          end
        end
      end else begin
        if(when_SuperResolutionPart3_l694) begin
          if(when_SuperResolutionPart3_l697) begin
            if(compareStage_controlPipe_payload_lastRow) begin
              if(compareStage_controlPipe_payload_counterCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_mainThreePixelStream_payload - compareStage_counterThreePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterThreePixelStream_payload - compareStage_mainThreePixelStream_payload);
              end
            end else begin
              if(compareStage_controlPipe_payload_counterCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_mainOnePixelStream_payload - compareStage_counterThreePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterThreePixelStream_payload - compareStage_mainOnePixelStream_payload);
              end
            end
          end else begin
            if(compareStage_controlPipe_payload_lastRow) begin
              if(compareStage_controlPipe_payload_counterCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_mainOnePixelStream_payload - compareStage_counterOnePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterOnePixelStream_payload - compareStage_mainOnePixelStream_payload);
              end
            end else begin
              if(compareStage_controlPipe_payload_counterCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_mainThreePixelStream_payload - compareStage_counterOnePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterOnePixelStream_payload - compareStage_mainThreePixelStream_payload);
              end
            end
          end
        end else begin
          if(when_SuperResolutionPart3_l725) begin
            if(compareStage_controlPipe_payload_lastRow) begin
              if(compareStage_controlPipe_payload_counterCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterTwoPixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainTwoPixelStream_payload);
              end
            end else begin
              if(compareStage_controlPipe_payload_counterCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_mainOnePixelStream_payload - compareStage_counterTwoPixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainOnePixelStream_payload);
              end
            end
          end else begin
            if(compareStage_controlPipe_payload_lastRow) begin
              if(compareStage_controlPipe_payload_counterCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_mainOnePixelStream_payload - compareStage_counterOnePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterOnePixelStream_payload - compareStage_mainOnePixelStream_payload);
              end
            end else begin
              if(compareStage_controlPipe_payload_counterCompare) begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterOnePixelStream_payload);
              end else begin
                CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterOnePixelStream_payload - compareStage_mainTwoPixelStream_payload);
              end
            end
          end
        end
      end
    end
  end

  always @(*) begin
    CICC1851_compareStage_controlPipe_translated_payload_horizontalDiff = compareStage_controlPipe_payload_horizontalDiff;
    if(!compareStage_controlPipe_payload_finalResult) begin
      if(when_SuperResolutionPart3_l661) begin
        if(compareStage_controlPipe_payload_horizontalCompare) begin
          CICC1851_compareStage_controlPipe_translated_payload_horizontalDiff = (compareStage_mainOnePixelStream_payload - compareStage_counterOnePixelStream_payload);
        end else begin
          CICC1851_compareStage_controlPipe_translated_payload_horizontalDiff = (compareStage_counterOnePixelStream_payload - compareStage_mainOnePixelStream_payload);
        end
      end else begin
        if(when_SuperResolutionPart3_l694) begin
          if(compareStage_controlPipe_payload_horizontalCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_horizontalDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterTwoPixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_horizontalDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainTwoPixelStream_payload);
          end
        end else begin
          if(compareStage_controlPipe_payload_horizontalCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_horizontalDiff = (compareStage_mainThreePixelStream_payload - compareStage_counterThreePixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_horizontalDiff = (compareStage_counterThreePixelStream_payload - compareStage_mainThreePixelStream_payload);
          end
        end
      end
    end
  end

  always @(*) begin
    CICC1851_compareStage_controlPipe_translated_payload_verticalDiff = compareStage_controlPipe_payload_verticalDiff;
    if(compareStage_controlPipe_payload_finalResult) begin
      if(when_SuperResolutionPart3_l647) begin
        CICC1851_compareStage_controlPipe_translated_payload_verticalDiff = 8'h0;
      end else begin
        if(when_SuperResolutionPart3_l649) begin
          if(compareStage_controlPipe_payload_verticalCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_verticalDiff = (compareStage_mainTwoPixelStream_payload - compareStage_mainThreePixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_verticalDiff = (compareStage_mainThreePixelStream_payload - compareStage_mainTwoPixelStream_payload);
          end
        end else begin
          if(when_SuperResolutionPart3_l652) begin
            if(compareStage_controlPipe_payload_verticalCompare) begin
              CICC1851_compareStage_controlPipe_translated_payload_verticalDiff = (compareStage_mainOnePixelStream_payload - compareStage_mainThreePixelStream_payload);
            end else begin
              CICC1851_compareStage_controlPipe_translated_payload_verticalDiff = (compareStage_mainThreePixelStream_payload - compareStage_mainOnePixelStream_payload);
            end
          end else begin
            if(compareStage_controlPipe_payload_verticalCompare) begin
              CICC1851_compareStage_controlPipe_translated_payload_verticalDiff = (compareStage_mainOnePixelStream_payload - compareStage_mainTwoPixelStream_payload);
            end else begin
              CICC1851_compareStage_controlPipe_translated_payload_verticalDiff = (compareStage_mainTwoPixelStream_payload - compareStage_mainOnePixelStream_payload);
            end
          end
        end
      end
    end
  end

  always @(*) begin
    CICC1851_compareStage_controlPipe_translated_payload_inValidMinDiff = compareStage_controlPipe_payload_inValidMinDiff;
    if(when_SuperResolutionPart3_l753) begin
      CICC1851_compareStage_controlPipe_translated_payload_inValidMinDiff = 1'b1;
    end
  end

  assign when_SuperResolutionPart3_l647 = (compareStage_controlPipe_payload_firstRow || compareStage_controlPipe_payload_lastRow);
  assign when_SuperResolutionPart3_l649 = (compareStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l652 = (compareStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l661 = (compareStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l664 = (compareStage_controlPipe_payload_nextPosition == 2'b01);
  assign when_SuperResolutionPart3_l697 = (compareStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l725 = (compareStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l694 = (compareStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l753 = ((((! compareStage_controlPipe_payload_finalResult) && (! compareStage_controlPipe_payload_mainDirectionValid)) && (! compareStage_controlPipe_payload_counterDirectionValid)) && (! compareStage_controlPipe_payload_horizontalDirectionValid));
  assign compareStage_controlPipe_translated_valid = compareStage_controlPipe_valid;
  assign compareStage_controlPipe_ready = compareStage_controlPipe_translated_ready;
  assign compareStage_controlPipe_translated_payload_frameStart = compareStage_controlPipe_payload_frameStart;
  assign compareStage_controlPipe_translated_payload_rowEnd = compareStage_controlPipe_payload_rowEnd;
  assign compareStage_controlPipe_translated_payload_pipeValid = compareStage_controlPipe_payload_pipeValid;
  assign compareStage_controlPipe_translated_payload_firstRow = compareStage_controlPipe_payload_firstRow;
  assign compareStage_controlPipe_translated_payload_lastRow = compareStage_controlPipe_payload_lastRow;
  assign compareStage_controlPipe_translated_payload_finalResult = compareStage_controlPipe_payload_finalResult;
  assign compareStage_controlPipe_translated_payload_mainCompare = compareStage_controlPipe_payload_mainCompare;
  assign compareStage_controlPipe_translated_payload_counterCompare = compareStage_controlPipe_payload_counterCompare;
  assign compareStage_controlPipe_translated_payload_horizontalCompare = compareStage_controlPipe_payload_horizontalCompare;
  assign compareStage_controlPipe_translated_payload_verticalCompare = compareStage_controlPipe_payload_verticalCompare;
  assign compareStage_controlPipe_translated_payload_mainDiff = CICC1851_compareStage_controlPipe_translated_payload_mainDiff;
  assign compareStage_controlPipe_translated_payload_counterDiff = CICC1851_compareStage_controlPipe_translated_payload_counterDiff;
  assign compareStage_controlPipe_translated_payload_horizontalDiff = CICC1851_compareStage_controlPipe_translated_payload_horizontalDiff;
  assign compareStage_controlPipe_translated_payload_verticalDiff = CICC1851_compareStage_controlPipe_translated_payload_verticalDiff;
  assign compareStage_controlPipe_translated_payload_isHorizontalMin = compareStage_controlPipe_payload_isHorizontalMin;
  assign compareStage_controlPipe_translated_payload_minDiff = compareStage_controlPipe_payload_minDiff;
  assign compareStage_controlPipe_translated_payload_currentPosition = compareStage_controlPipe_payload_currentPosition;
  assign compareStage_controlPipe_translated_payload_nextPosition = compareStage_controlPipe_payload_nextPosition;
  assign compareStage_controlPipe_translated_payload_horizontalDirectionValid = compareStage_controlPipe_payload_horizontalDirectionValid;
  assign compareStage_controlPipe_translated_payload_verticalDirectionValid = compareStage_controlPipe_payload_verticalDirectionValid;
  assign compareStage_controlPipe_translated_payload_mainDirectionValid = compareStage_controlPipe_payload_mainDirectionValid;
  assign compareStage_controlPipe_translated_payload_counterDirectionValid = compareStage_controlPipe_payload_counterDirectionValid;
  assign compareStage_controlPipe_translated_payload_inValidMinDiff = CICC1851_compareStage_controlPipe_translated_payload_inValidMinDiff;
  assign compareStage_controlPipe_translated_ready = (! compareStage_controlPipe_translated_rValid);
  assign compareStage_controlPipe_translated_s2mPipe_valid = (compareStage_controlPipe_translated_valid || compareStage_controlPipe_translated_rValid);
  assign compareStage_controlPipe_translated_s2mPipe_payload_frameStart = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_frameStart : compareStage_controlPipe_translated_payload_frameStart);
  assign compareStage_controlPipe_translated_s2mPipe_payload_rowEnd = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_rowEnd : compareStage_controlPipe_translated_payload_rowEnd);
  assign compareStage_controlPipe_translated_s2mPipe_payload_pipeValid = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_pipeValid : compareStage_controlPipe_translated_payload_pipeValid);
  assign compareStage_controlPipe_translated_s2mPipe_payload_firstRow = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_firstRow : compareStage_controlPipe_translated_payload_firstRow);
  assign compareStage_controlPipe_translated_s2mPipe_payload_lastRow = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_lastRow : compareStage_controlPipe_translated_payload_lastRow);
  assign compareStage_controlPipe_translated_s2mPipe_payload_finalResult = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_finalResult : compareStage_controlPipe_translated_payload_finalResult);
  assign compareStage_controlPipe_translated_s2mPipe_payload_mainCompare = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_mainCompare : compareStage_controlPipe_translated_payload_mainCompare);
  assign compareStage_controlPipe_translated_s2mPipe_payload_counterCompare = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_counterCompare : compareStage_controlPipe_translated_payload_counterCompare);
  assign compareStage_controlPipe_translated_s2mPipe_payload_horizontalCompare = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_horizontalCompare : compareStage_controlPipe_translated_payload_horizontalCompare);
  assign compareStage_controlPipe_translated_s2mPipe_payload_verticalCompare = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_verticalCompare : compareStage_controlPipe_translated_payload_verticalCompare);
  assign compareStage_controlPipe_translated_s2mPipe_payload_mainDiff = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_mainDiff : compareStage_controlPipe_translated_payload_mainDiff);
  assign compareStage_controlPipe_translated_s2mPipe_payload_counterDiff = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_counterDiff : compareStage_controlPipe_translated_payload_counterDiff);
  assign compareStage_controlPipe_translated_s2mPipe_payload_horizontalDiff = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_horizontalDiff : compareStage_controlPipe_translated_payload_horizontalDiff);
  assign compareStage_controlPipe_translated_s2mPipe_payload_verticalDiff = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_verticalDiff : compareStage_controlPipe_translated_payload_verticalDiff);
  assign compareStage_controlPipe_translated_s2mPipe_payload_isHorizontalMin = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_isHorizontalMin : compareStage_controlPipe_translated_payload_isHorizontalMin);
  assign compareStage_controlPipe_translated_s2mPipe_payload_minDiff = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_minDiff : compareStage_controlPipe_translated_payload_minDiff);
  assign compareStage_controlPipe_translated_s2mPipe_payload_currentPosition = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_currentPosition : compareStage_controlPipe_translated_payload_currentPosition);
  assign compareStage_controlPipe_translated_s2mPipe_payload_nextPosition = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_nextPosition : compareStage_controlPipe_translated_payload_nextPosition);
  assign compareStage_controlPipe_translated_s2mPipe_payload_horizontalDirectionValid = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_horizontalDirectionValid : compareStage_controlPipe_translated_payload_horizontalDirectionValid);
  assign compareStage_controlPipe_translated_s2mPipe_payload_verticalDirectionValid = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_verticalDirectionValid : compareStage_controlPipe_translated_payload_verticalDirectionValid);
  assign compareStage_controlPipe_translated_s2mPipe_payload_mainDirectionValid = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_mainDirectionValid : compareStage_controlPipe_translated_payload_mainDirectionValid);
  assign compareStage_controlPipe_translated_s2mPipe_payload_counterDirectionValid = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_counterDirectionValid : compareStage_controlPipe_translated_payload_counterDirectionValid);
  assign compareStage_controlPipe_translated_s2mPipe_payload_inValidMinDiff = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_inValidMinDiff : compareStage_controlPipe_translated_payload_inValidMinDiff);
  always @(*) begin
    compareStage_controlPipe_translated_s2mPipe_ready = diffStage_controlPipe_ready;
    if(when_Stream_l368_53) begin
      compareStage_controlPipe_translated_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_53 = (! diffStage_controlPipe_valid);
  assign diffStage_controlPipe_valid = compareStage_controlPipe_translated_s2mPipe_rValid;
  assign diffStage_controlPipe_payload_frameStart = compareStage_controlPipe_translated_s2mPipe_rData_frameStart;
  assign diffStage_controlPipe_payload_rowEnd = compareStage_controlPipe_translated_s2mPipe_rData_rowEnd;
  assign diffStage_controlPipe_payload_pipeValid = compareStage_controlPipe_translated_s2mPipe_rData_pipeValid;
  assign diffStage_controlPipe_payload_firstRow = compareStage_controlPipe_translated_s2mPipe_rData_firstRow;
  assign diffStage_controlPipe_payload_lastRow = compareStage_controlPipe_translated_s2mPipe_rData_lastRow;
  assign diffStage_controlPipe_payload_finalResult = compareStage_controlPipe_translated_s2mPipe_rData_finalResult;
  assign diffStage_controlPipe_payload_mainCompare = compareStage_controlPipe_translated_s2mPipe_rData_mainCompare;
  assign diffStage_controlPipe_payload_counterCompare = compareStage_controlPipe_translated_s2mPipe_rData_counterCompare;
  assign diffStage_controlPipe_payload_horizontalCompare = compareStage_controlPipe_translated_s2mPipe_rData_horizontalCompare;
  assign diffStage_controlPipe_payload_verticalCompare = compareStage_controlPipe_translated_s2mPipe_rData_verticalCompare;
  assign diffStage_controlPipe_payload_mainDiff = compareStage_controlPipe_translated_s2mPipe_rData_mainDiff;
  assign diffStage_controlPipe_payload_counterDiff = compareStage_controlPipe_translated_s2mPipe_rData_counterDiff;
  assign diffStage_controlPipe_payload_horizontalDiff = compareStage_controlPipe_translated_s2mPipe_rData_horizontalDiff;
  assign diffStage_controlPipe_payload_verticalDiff = compareStage_controlPipe_translated_s2mPipe_rData_verticalDiff;
  assign diffStage_controlPipe_payload_isHorizontalMin = compareStage_controlPipe_translated_s2mPipe_rData_isHorizontalMin;
  assign diffStage_controlPipe_payload_minDiff = compareStage_controlPipe_translated_s2mPipe_rData_minDiff;
  assign diffStage_controlPipe_payload_currentPosition = compareStage_controlPipe_translated_s2mPipe_rData_currentPosition;
  assign diffStage_controlPipe_payload_nextPosition = compareStage_controlPipe_translated_s2mPipe_rData_nextPosition;
  assign diffStage_controlPipe_payload_horizontalDirectionValid = compareStage_controlPipe_translated_s2mPipe_rData_horizontalDirectionValid;
  assign diffStage_controlPipe_payload_verticalDirectionValid = compareStage_controlPipe_translated_s2mPipe_rData_verticalDirectionValid;
  assign diffStage_controlPipe_payload_mainDirectionValid = compareStage_controlPipe_translated_s2mPipe_rData_mainDirectionValid;
  assign diffStage_controlPipe_payload_counterDirectionValid = compareStage_controlPipe_translated_s2mPipe_rData_counterDirectionValid;
  assign diffStage_controlPipe_payload_inValidMinDiff = compareStage_controlPipe_translated_s2mPipe_rData_inValidMinDiff;
  assign diffStage_mainOnePixelStream_ready = (! diffStage_mainOnePixelStream_rValid);
  assign diffStage_mainOnePixelStream_s2mPipe_valid = (diffStage_mainOnePixelStream_valid || diffStage_mainOnePixelStream_rValid);
  assign diffStage_mainOnePixelStream_s2mPipe_payload = (diffStage_mainOnePixelStream_rValid ? diffStage_mainOnePixelStream_rData : diffStage_mainOnePixelStream_payload);
  always @(*) begin
    diffStage_mainOnePixelStream_s2mPipe_ready = resultStage_mainOnePixelStream_ready;
    if(when_Stream_l368_54) begin
      diffStage_mainOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_54 = (! resultStage_mainOnePixelStream_valid);
  assign resultStage_mainOnePixelStream_valid = diffStage_mainOnePixelStream_s2mPipe_rValid;
  assign resultStage_mainOnePixelStream_payload = diffStage_mainOnePixelStream_s2mPipe_rData;
  assign diffStage_counterOnePixelStream_ready = (! diffStage_counterOnePixelStream_rValid);
  assign diffStage_counterOnePixelStream_s2mPipe_valid = (diffStage_counterOnePixelStream_valid || diffStage_counterOnePixelStream_rValid);
  assign diffStage_counterOnePixelStream_s2mPipe_payload = (diffStage_counterOnePixelStream_rValid ? diffStage_counterOnePixelStream_rData : diffStage_counterOnePixelStream_payload);
  always @(*) begin
    diffStage_counterOnePixelStream_s2mPipe_ready = resultStage_counterOnePixelStream_ready;
    if(when_Stream_l368_55) begin
      diffStage_counterOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_55 = (! resultStage_counterOnePixelStream_valid);
  assign resultStage_counterOnePixelStream_valid = diffStage_counterOnePixelStream_s2mPipe_rValid;
  assign resultStage_counterOnePixelStream_payload = diffStage_counterOnePixelStream_s2mPipe_rData;
  assign diffStage_mainTwoPixelStream_ready = (! diffStage_mainTwoPixelStream_rValid);
  assign diffStage_mainTwoPixelStream_s2mPipe_valid = (diffStage_mainTwoPixelStream_valid || diffStage_mainTwoPixelStream_rValid);
  assign diffStage_mainTwoPixelStream_s2mPipe_payload = (diffStage_mainTwoPixelStream_rValid ? diffStage_mainTwoPixelStream_rData : diffStage_mainTwoPixelStream_payload);
  always @(*) begin
    diffStage_mainTwoPixelStream_s2mPipe_ready = resultStage_mainTwoPixelStream_ready;
    if(when_Stream_l368_56) begin
      diffStage_mainTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_56 = (! resultStage_mainTwoPixelStream_valid);
  assign resultStage_mainTwoPixelStream_valid = diffStage_mainTwoPixelStream_s2mPipe_rValid;
  assign resultStage_mainTwoPixelStream_payload = diffStage_mainTwoPixelStream_s2mPipe_rData;
  assign diffStage_counterTwoPixelStream_ready = (! diffStage_counterTwoPixelStream_rValid);
  assign diffStage_counterTwoPixelStream_s2mPipe_valid = (diffStage_counterTwoPixelStream_valid || diffStage_counterTwoPixelStream_rValid);
  assign diffStage_counterTwoPixelStream_s2mPipe_payload = (diffStage_counterTwoPixelStream_rValid ? diffStage_counterTwoPixelStream_rData : diffStage_counterTwoPixelStream_payload);
  always @(*) begin
    diffStage_counterTwoPixelStream_s2mPipe_ready = resultStage_counterTwoPixelStream_ready;
    if(when_Stream_l368_57) begin
      diffStage_counterTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_57 = (! resultStage_counterTwoPixelStream_valid);
  assign resultStage_counterTwoPixelStream_valid = diffStage_counterTwoPixelStream_s2mPipe_rValid;
  assign resultStage_counterTwoPixelStream_payload = diffStage_counterTwoPixelStream_s2mPipe_rData;
  assign diffStage_mainThreePixelStream_ready = (! diffStage_mainThreePixelStream_rValid);
  assign diffStage_mainThreePixelStream_s2mPipe_valid = (diffStage_mainThreePixelStream_valid || diffStage_mainThreePixelStream_rValid);
  assign diffStage_mainThreePixelStream_s2mPipe_payload = (diffStage_mainThreePixelStream_rValid ? diffStage_mainThreePixelStream_rData : diffStage_mainThreePixelStream_payload);
  always @(*) begin
    diffStage_mainThreePixelStream_s2mPipe_ready = resultStage_mainThreePixelStream_ready;
    if(when_Stream_l368_58) begin
      diffStage_mainThreePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_58 = (! resultStage_mainThreePixelStream_valid);
  assign resultStage_mainThreePixelStream_valid = diffStage_mainThreePixelStream_s2mPipe_rValid;
  assign resultStage_mainThreePixelStream_payload = diffStage_mainThreePixelStream_s2mPipe_rData;
  assign diffStage_counterThreePixelStream_ready = (! diffStage_counterThreePixelStream_rValid);
  assign diffStage_counterThreePixelStream_s2mPipe_valid = (diffStage_counterThreePixelStream_valid || diffStage_counterThreePixelStream_rValid);
  assign diffStage_counterThreePixelStream_s2mPipe_payload = (diffStage_counterThreePixelStream_rValid ? diffStage_counterThreePixelStream_rData : diffStage_counterThreePixelStream_payload);
  always @(*) begin
    diffStage_counterThreePixelStream_s2mPipe_ready = resultStage_counterThreePixelStream_ready;
    if(when_Stream_l368_59) begin
      diffStage_counterThreePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_59 = (! resultStage_counterThreePixelStream_valid);
  assign resultStage_counterThreePixelStream_valid = diffStage_counterThreePixelStream_s2mPipe_rValid;
  assign resultStage_counterThreePixelStream_payload = diffStage_counterThreePixelStream_s2mPipe_rData;
  assign diffStage_mainOneValidStream_ready = (! diffStage_mainOneValidStream_rValid);
  assign diffStage_mainOneValidStream_s2mPipe_valid = (diffStage_mainOneValidStream_valid || diffStage_mainOneValidStream_rValid);
  assign diffStage_mainOneValidStream_s2mPipe_payload = (diffStage_mainOneValidStream_rValid ? diffStage_mainOneValidStream_rData : diffStage_mainOneValidStream_payload);
  always @(*) begin
    diffStage_mainOneValidStream_s2mPipe_ready = resultStage_mainOneValidStream_ready;
    if(when_Stream_l368_60) begin
      diffStage_mainOneValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_60 = (! resultStage_mainOneValidStream_valid);
  assign resultStage_mainOneValidStream_valid = diffStage_mainOneValidStream_s2mPipe_rValid;
  assign resultStage_mainOneValidStream_payload = diffStage_mainOneValidStream_s2mPipe_rData;
  assign diffStage_counterOneValidStream_ready = (! diffStage_counterOneValidStream_rValid);
  assign diffStage_counterOneValidStream_s2mPipe_valid = (diffStage_counterOneValidStream_valid || diffStage_counterOneValidStream_rValid);
  assign diffStage_counterOneValidStream_s2mPipe_payload = (diffStage_counterOneValidStream_rValid ? diffStage_counterOneValidStream_rData : diffStage_counterOneValidStream_payload);
  always @(*) begin
    diffStage_counterOneValidStream_s2mPipe_ready = resultStage_counterOneValidStream_ready;
    if(when_Stream_l368_61) begin
      diffStage_counterOneValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_61 = (! resultStage_counterOneValidStream_valid);
  assign resultStage_counterOneValidStream_valid = diffStage_counterOneValidStream_s2mPipe_rValid;
  assign resultStage_counterOneValidStream_payload = diffStage_counterOneValidStream_s2mPipe_rData;
  assign diffStage_mainTwoValidStream_ready = (! diffStage_mainTwoValidStream_rValid);
  assign diffStage_mainTwoValidStream_s2mPipe_valid = (diffStage_mainTwoValidStream_valid || diffStage_mainTwoValidStream_rValid);
  assign diffStage_mainTwoValidStream_s2mPipe_payload = (diffStage_mainTwoValidStream_rValid ? diffStage_mainTwoValidStream_rData : diffStage_mainTwoValidStream_payload);
  always @(*) begin
    diffStage_mainTwoValidStream_s2mPipe_ready = resultStage_mainTwoValidStream_ready;
    if(when_Stream_l368_62) begin
      diffStage_mainTwoValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_62 = (! resultStage_mainTwoValidStream_valid);
  assign resultStage_mainTwoValidStream_valid = diffStage_mainTwoValidStream_s2mPipe_rValid;
  assign resultStage_mainTwoValidStream_payload = diffStage_mainTwoValidStream_s2mPipe_rData;
  assign diffStage_counterTwoValidStream_ready = (! diffStage_counterTwoValidStream_rValid);
  assign diffStage_counterTwoValidStream_s2mPipe_valid = (diffStage_counterTwoValidStream_valid || diffStage_counterTwoValidStream_rValid);
  assign diffStage_counterTwoValidStream_s2mPipe_payload = (diffStage_counterTwoValidStream_rValid ? diffStage_counterTwoValidStream_rData : diffStage_counterTwoValidStream_payload);
  always @(*) begin
    diffStage_counterTwoValidStream_s2mPipe_ready = resultStage_counterTwoValidStream_ready;
    if(when_Stream_l368_63) begin
      diffStage_counterTwoValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_63 = (! resultStage_counterTwoValidStream_valid);
  assign resultStage_counterTwoValidStream_valid = diffStage_counterTwoValidStream_s2mPipe_rValid;
  assign resultStage_counterTwoValidStream_payload = diffStage_counterTwoValidStream_s2mPipe_rData;
  assign diffStage_mainThreeValidStream_ready = (! diffStage_mainThreeValidStream_rValid);
  assign diffStage_mainThreeValidStream_s2mPipe_valid = (diffStage_mainThreeValidStream_valid || diffStage_mainThreeValidStream_rValid);
  assign diffStage_mainThreeValidStream_s2mPipe_payload = (diffStage_mainThreeValidStream_rValid ? diffStage_mainThreeValidStream_rData : diffStage_mainThreeValidStream_payload);
  always @(*) begin
    diffStage_mainThreeValidStream_s2mPipe_ready = resultStage_mainThreeValidStream_ready;
    if(when_Stream_l368_64) begin
      diffStage_mainThreeValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_64 = (! resultStage_mainThreeValidStream_valid);
  assign resultStage_mainThreeValidStream_valid = diffStage_mainThreeValidStream_s2mPipe_rValid;
  assign resultStage_mainThreeValidStream_payload = diffStage_mainThreeValidStream_s2mPipe_rData;
  assign diffStage_counterThreeValidStream_ready = (! diffStage_counterThreeValidStream_rValid);
  assign diffStage_counterThreeValidStream_s2mPipe_valid = (diffStage_counterThreeValidStream_valid || diffStage_counterThreeValidStream_rValid);
  assign diffStage_counterThreeValidStream_s2mPipe_payload = (diffStage_counterThreeValidStream_rValid ? diffStage_counterThreeValidStream_rData : diffStage_counterThreeValidStream_payload);
  always @(*) begin
    diffStage_counterThreeValidStream_s2mPipe_ready = resultStage_counterThreeValidStream_ready;
    if(when_Stream_l368_65) begin
      diffStage_counterThreeValidStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_65 = (! resultStage_counterThreeValidStream_valid);
  assign resultStage_counterThreeValidStream_valid = diffStage_counterThreeValidStream_s2mPipe_rValid;
  assign resultStage_counterThreeValidStream_payload = diffStage_counterThreeValidStream_s2mPipe_rData;
  assign diffStage_controlPipe_ready = diffStage_controlPipe_fork_io_input_ready;
  always @(*) begin
    CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin = diffStage_controlPipe_payload_isHorizontalMin;
    if(when_SuperResolutionPart3_l783) begin
      if(when_SuperResolutionPart3_l784) begin
        if(when_SuperResolutionPart3_l785) begin
          CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin = 1'b1;
        end else begin
          if(when_SuperResolutionPart3_l788) begin
            CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin = 1'b0;
          end else begin
            CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin = 1'b0;
          end
        end
      end else begin
        if(when_SuperResolutionPart3_l795) begin
          if(when_SuperResolutionPart3_l796) begin
            CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin = 1'b0;
          end else begin
            CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin = 1'b0;
          end
        end else begin
          if(when_SuperResolutionPart3_l803) begin
            if(when_SuperResolutionPart3_l804) begin
              CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin = 1'b1;
            end else begin
              CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin = 1'b0;
            end
          end else begin
            if(when_SuperResolutionPart3_l811) begin
              if(when_SuperResolutionPart3_l812) begin
                CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin = 1'b1;
              end else begin
                CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin = 1'b0;
              end
            end else begin
              if(when_SuperResolutionPart3_l819) begin
                CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin = 1'b0;
              end else begin
                if(when_SuperResolutionPart3_l822) begin
                  CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin = 1'b1;
                end else begin
                  if(when_SuperResolutionPart3_l825) begin
                    CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin = 1'b0;
                  end
                end
              end
            end
          end
        end
      end
    end
  end

  always @(*) begin
    CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff = diffStage_controlPipe_payload_minDiff;
    if(when_SuperResolutionPart3_l783) begin
      if(when_SuperResolutionPart3_l784) begin
        if(when_SuperResolutionPart3_l785) begin
          CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff = diffStage_controlPipe_payload_horizontalDiff;
        end else begin
          if(when_SuperResolutionPart3_l788) begin
            CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff = diffStage_controlPipe_payload_mainDiff;
          end else begin
            CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff = diffStage_controlPipe_payload_counterDiff;
          end
        end
      end else begin
        if(when_SuperResolutionPart3_l795) begin
          if(when_SuperResolutionPart3_l796) begin
            CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff = diffStage_controlPipe_payload_mainDiff;
          end else begin
            CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff = diffStage_controlPipe_payload_counterDiff;
          end
        end else begin
          if(when_SuperResolutionPart3_l803) begin
            if(when_SuperResolutionPart3_l804) begin
              CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff = diffStage_controlPipe_payload_horizontalDiff;
            end else begin
              CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff = diffStage_controlPipe_payload_counterDiff;
            end
          end else begin
            if(when_SuperResolutionPart3_l811) begin
              if(when_SuperResolutionPart3_l812) begin
                CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff = diffStage_controlPipe_payload_horizontalDiff;
              end else begin
                CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff = diffStage_controlPipe_payload_mainDiff;
              end
            end else begin
              if(when_SuperResolutionPart3_l819) begin
                CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff = diffStage_controlPipe_payload_counterDiff;
              end else begin
                if(when_SuperResolutionPart3_l822) begin
                  CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff = diffStage_controlPipe_payload_horizontalDiff;
                end else begin
                  if(when_SuperResolutionPart3_l825) begin
                    CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff = diffStage_controlPipe_payload_mainDiff;
                  end
                end
              end
            end
          end
        end
      end
    end
  end

  assign when_SuperResolutionPart3_l783 = (! diffStage_controlPipe_payload_finalResult);
  assign when_SuperResolutionPart3_l784 = ((diffStage_controlPipe_payload_horizontalDirectionValid && diffStage_controlPipe_payload_mainDirectionValid) && diffStage_controlPipe_payload_counterDirectionValid);
  assign when_SuperResolutionPart3_l785 = ((diffStage_controlPipe_payload_horizontalDiff <= diffStage_controlPipe_payload_mainDiff) && (diffStage_controlPipe_payload_horizontalDiff <= diffStage_controlPipe_payload_counterDiff));
  assign when_SuperResolutionPart3_l788 = ((diffStage_controlPipe_payload_mainDiff < diffStage_controlPipe_payload_horizontalDiff) && (diffStage_controlPipe_payload_mainDiff <= diffStage_controlPipe_payload_counterDiff));
  assign when_SuperResolutionPart3_l796 = (diffStage_controlPipe_payload_mainDiff <= diffStage_controlPipe_payload_counterDiff);
  assign when_SuperResolutionPart3_l804 = (diffStage_controlPipe_payload_horizontalDiff <= diffStage_controlPipe_payload_counterDiff);
  assign when_SuperResolutionPart3_l812 = (diffStage_controlPipe_payload_horizontalDiff <= diffStage_controlPipe_payload_mainDiff);
  assign when_SuperResolutionPart3_l795 = (((! diffStage_controlPipe_payload_horizontalDirectionValid) && diffStage_controlPipe_payload_mainDirectionValid) && diffStage_controlPipe_payload_counterDirectionValid);
  assign when_SuperResolutionPart3_l803 = ((diffStage_controlPipe_payload_horizontalDirectionValid && (! diffStage_controlPipe_payload_mainDirectionValid)) && diffStage_controlPipe_payload_counterDirectionValid);
  assign when_SuperResolutionPart3_l811 = ((diffStage_controlPipe_payload_horizontalDirectionValid && diffStage_controlPipe_payload_mainDirectionValid) && (! diffStage_controlPipe_payload_counterDirectionValid));
  assign when_SuperResolutionPart3_l819 = (((! diffStage_controlPipe_payload_horizontalDirectionValid) && (! diffStage_controlPipe_payload_mainDirectionValid)) && diffStage_controlPipe_payload_counterDirectionValid);
  assign when_SuperResolutionPart3_l822 = ((diffStage_controlPipe_payload_horizontalDirectionValid && (! diffStage_controlPipe_payload_mainDirectionValid)) && (! diffStage_controlPipe_payload_counterDirectionValid));
  assign when_SuperResolutionPart3_l825 = (((! diffStage_controlPipe_payload_horizontalDirectionValid) && diffStage_controlPipe_payload_mainDirectionValid) && (! diffStage_controlPipe_payload_counterDirectionValid));
  assign resultStage_controlPipeBeforePipe_valid = diffStage_controlPipe_fork_io_outputs_0_valid;
  assign resultStage_controlPipeBeforePipe_payload_frameStart = diffStage_controlPipe_payload_frameStart;
  assign resultStage_controlPipeBeforePipe_payload_rowEnd = diffStage_controlPipe_payload_rowEnd;
  assign resultStage_controlPipeBeforePipe_payload_pipeValid = diffStage_controlPipe_payload_pipeValid;
  assign resultStage_controlPipeBeforePipe_payload_firstRow = diffStage_controlPipe_payload_firstRow;
  assign resultStage_controlPipeBeforePipe_payload_lastRow = diffStage_controlPipe_payload_lastRow;
  assign resultStage_controlPipeBeforePipe_payload_finalResult = diffStage_controlPipe_payload_finalResult;
  assign resultStage_controlPipeBeforePipe_payload_mainCompare = diffStage_controlPipe_payload_mainCompare;
  assign resultStage_controlPipeBeforePipe_payload_counterCompare = diffStage_controlPipe_payload_counterCompare;
  assign resultStage_controlPipeBeforePipe_payload_horizontalCompare = diffStage_controlPipe_payload_horizontalCompare;
  assign resultStage_controlPipeBeforePipe_payload_verticalCompare = diffStage_controlPipe_payload_verticalCompare;
  assign resultStage_controlPipeBeforePipe_payload_mainDiff = diffStage_controlPipe_payload_mainDiff;
  assign resultStage_controlPipeBeforePipe_payload_counterDiff = diffStage_controlPipe_payload_counterDiff;
  assign resultStage_controlPipeBeforePipe_payload_horizontalDiff = diffStage_controlPipe_payload_horizontalDiff;
  assign resultStage_controlPipeBeforePipe_payload_verticalDiff = diffStage_controlPipe_payload_verticalDiff;
  assign resultStage_controlPipeBeforePipe_payload_isHorizontalMin = CICC1851_resultStage_controlPipeBeforePipe_payload_isHorizontalMin;
  assign resultStage_controlPipeBeforePipe_payload_minDiff = CICC1851_resultStage_controlPipeBeforePipe_payload_minDiff;
  assign resultStage_controlPipeBeforePipe_payload_currentPosition = diffStage_controlPipe_payload_currentPosition;
  assign resultStage_controlPipeBeforePipe_payload_nextPosition = diffStage_controlPipe_payload_nextPosition;
  assign resultStage_controlPipeBeforePipe_payload_horizontalDirectionValid = diffStage_controlPipe_payload_horizontalDirectionValid;
  assign resultStage_controlPipeBeforePipe_payload_verticalDirectionValid = diffStage_controlPipe_payload_verticalDirectionValid;
  assign resultStage_controlPipeBeforePipe_payload_mainDirectionValid = diffStage_controlPipe_payload_mainDirectionValid;
  assign resultStage_controlPipeBeforePipe_payload_counterDirectionValid = diffStage_controlPipe_payload_counterDirectionValid;
  assign resultStage_controlPipeBeforePipe_payload_inValidMinDiff = diffStage_controlPipe_payload_inValidMinDiff;
  assign resultStage_controlPipeBeforePipe_ready = (! resultStage_controlPipeBeforePipe_rValid);
  assign resultStage_controlPipeBeforePipe_s2mPipe_valid = (resultStage_controlPipeBeforePipe_valid || resultStage_controlPipeBeforePipe_rValid);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_frameStart = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_frameStart : resultStage_controlPipeBeforePipe_payload_frameStart);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_rowEnd = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_rowEnd : resultStage_controlPipeBeforePipe_payload_rowEnd);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_pipeValid = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_pipeValid : resultStage_controlPipeBeforePipe_payload_pipeValid);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_firstRow = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_firstRow : resultStage_controlPipeBeforePipe_payload_firstRow);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_lastRow = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_lastRow : resultStage_controlPipeBeforePipe_payload_lastRow);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_finalResult = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_finalResult : resultStage_controlPipeBeforePipe_payload_finalResult);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_mainCompare = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_mainCompare : resultStage_controlPipeBeforePipe_payload_mainCompare);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_counterCompare = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_counterCompare : resultStage_controlPipeBeforePipe_payload_counterCompare);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_horizontalCompare = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_horizontalCompare : resultStage_controlPipeBeforePipe_payload_horizontalCompare);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_verticalCompare = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_verticalCompare : resultStage_controlPipeBeforePipe_payload_verticalCompare);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_mainDiff = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_mainDiff : resultStage_controlPipeBeforePipe_payload_mainDiff);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_counterDiff = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_counterDiff : resultStage_controlPipeBeforePipe_payload_counterDiff);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_horizontalDiff = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_horizontalDiff : resultStage_controlPipeBeforePipe_payload_horizontalDiff);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_verticalDiff = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_verticalDiff : resultStage_controlPipeBeforePipe_payload_verticalDiff);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_isHorizontalMin = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_isHorizontalMin : resultStage_controlPipeBeforePipe_payload_isHorizontalMin);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_minDiff = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_minDiff : resultStage_controlPipeBeforePipe_payload_minDiff);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_currentPosition = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_currentPosition : resultStage_controlPipeBeforePipe_payload_currentPosition);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_nextPosition = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_nextPosition : resultStage_controlPipeBeforePipe_payload_nextPosition);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_horizontalDirectionValid = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_horizontalDirectionValid : resultStage_controlPipeBeforePipe_payload_horizontalDirectionValid);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_verticalDirectionValid = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_verticalDirectionValid : resultStage_controlPipeBeforePipe_payload_verticalDirectionValid);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_mainDirectionValid = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_mainDirectionValid : resultStage_controlPipeBeforePipe_payload_mainDirectionValid);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_counterDirectionValid = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_counterDirectionValid : resultStage_controlPipeBeforePipe_payload_counterDirectionValid);
  assign resultStage_controlPipeBeforePipe_s2mPipe_payload_inValidMinDiff = (resultStage_controlPipeBeforePipe_rValid ? resultStage_controlPipeBeforePipe_rData_inValidMinDiff : resultStage_controlPipeBeforePipe_payload_inValidMinDiff);
  always @(*) begin
    resultStage_controlPipeBeforePipe_s2mPipe_ready = resultStage_controlPipe_ready;
    if(when_Stream_l368_66) begin
      resultStage_controlPipeBeforePipe_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_66 = (! resultStage_controlPipe_valid);
  assign resultStage_controlPipe_valid = resultStage_controlPipeBeforePipe_s2mPipe_rValid;
  assign resultStage_controlPipe_payload_frameStart = resultStage_controlPipeBeforePipe_s2mPipe_rData_frameStart;
  assign resultStage_controlPipe_payload_rowEnd = resultStage_controlPipeBeforePipe_s2mPipe_rData_rowEnd;
  assign resultStage_controlPipe_payload_pipeValid = resultStage_controlPipeBeforePipe_s2mPipe_rData_pipeValid;
  assign resultStage_controlPipe_payload_firstRow = resultStage_controlPipeBeforePipe_s2mPipe_rData_firstRow;
  assign resultStage_controlPipe_payload_lastRow = resultStage_controlPipeBeforePipe_s2mPipe_rData_lastRow;
  assign resultStage_controlPipe_payload_finalResult = resultStage_controlPipeBeforePipe_s2mPipe_rData_finalResult;
  assign resultStage_controlPipe_payload_mainCompare = resultStage_controlPipeBeforePipe_s2mPipe_rData_mainCompare;
  assign resultStage_controlPipe_payload_counterCompare = resultStage_controlPipeBeforePipe_s2mPipe_rData_counterCompare;
  assign resultStage_controlPipe_payload_horizontalCompare = resultStage_controlPipeBeforePipe_s2mPipe_rData_horizontalCompare;
  assign resultStage_controlPipe_payload_verticalCompare = resultStage_controlPipeBeforePipe_s2mPipe_rData_verticalCompare;
  assign resultStage_controlPipe_payload_mainDiff = resultStage_controlPipeBeforePipe_s2mPipe_rData_mainDiff;
  assign resultStage_controlPipe_payload_counterDiff = resultStage_controlPipeBeforePipe_s2mPipe_rData_counterDiff;
  assign resultStage_controlPipe_payload_horizontalDiff = resultStage_controlPipeBeforePipe_s2mPipe_rData_horizontalDiff;
  assign resultStage_controlPipe_payload_verticalDiff = resultStage_controlPipeBeforePipe_s2mPipe_rData_verticalDiff;
  assign resultStage_controlPipe_payload_isHorizontalMin = resultStage_controlPipeBeforePipe_s2mPipe_rData_isHorizontalMin;
  assign resultStage_controlPipe_payload_minDiff = resultStage_controlPipeBeforePipe_s2mPipe_rData_minDiff;
  assign resultStage_controlPipe_payload_currentPosition = resultStage_controlPipeBeforePipe_s2mPipe_rData_currentPosition;
  assign resultStage_controlPipe_payload_nextPosition = resultStage_controlPipeBeforePipe_s2mPipe_rData_nextPosition;
  assign resultStage_controlPipe_payload_horizontalDirectionValid = resultStage_controlPipeBeforePipe_s2mPipe_rData_horizontalDirectionValid;
  assign resultStage_controlPipe_payload_verticalDirectionValid = resultStage_controlPipeBeforePipe_s2mPipe_rData_verticalDirectionValid;
  assign resultStage_controlPipe_payload_mainDirectionValid = resultStage_controlPipeBeforePipe_s2mPipe_rData_mainDirectionValid;
  assign resultStage_controlPipe_payload_counterDirectionValid = resultStage_controlPipeBeforePipe_s2mPipe_rData_counterDirectionValid;
  assign resultStage_controlPipe_payload_inValidMinDiff = resultStage_controlPipeBeforePipe_s2mPipe_rData_inValidMinDiff;
  assign resultStage_pixelStream_valid = diffStage_controlPipe_fork_io_outputs_1_valid;
  always @(*) begin
    resultStage_pixelStream_payload = 8'h0;
    if(diffStage_controlPipe_payload_finalResult) begin
      if(when_SuperResolutionPart3_l840) begin
        resultStage_pixelStream_payload = diffStage_mainOnePixelStream_payload;
      end else begin
        if(when_SuperResolutionPart3_l841) begin
          resultStage_pixelStream_payload = diffStage_mainTwoPixelStream_payload;
        end else begin
          if(when_SuperResolutionPart3_l842) begin
            resultStage_pixelStream_payload = diffStage_mainThreePixelStream_payload;
          end else begin
            if(diffStage_controlPipe_payload_verticalDirectionValid) begin
              if(inValidMinDiff) begin
                if(when_SuperResolutionPart3_l846) begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload[7:0];
                end else begin
                  if(when_SuperResolutionPart3_l847) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_2[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_4[7:0];
                  end
                end
              end else begin
                if(when_SuperResolutionPart3_l850) begin
                  resultStage_pixelStream_payload = candidatePixel;
                end else begin
                  if(when_SuperResolutionPart3_l851) begin
                    if(isHorizontalDirection) begin
                      resultStage_pixelStream_payload = candidatePixel;
                    end else begin
                      if(when_SuperResolutionPart3_l854) begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_6[7:0];
                      end else begin
                        if(when_SuperResolutionPart3_l855) begin
                          resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_8[7:0];
                        end else begin
                          resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_10[7:0];
                        end
                      end
                    end
                  end else begin
                    if(when_SuperResolutionPart3_l860) begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_12[7:0];
                    end else begin
                      if(when_SuperResolutionPart3_l861) begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_14[7:0];
                      end else begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_16[7:0];
                      end
                    end
                  end
                end
              end
            end else begin
              resultStage_pixelStream_payload = candidatePixel;
            end
          end
        end
      end
    end else begin
      if(when_SuperResolutionPart3_l869) begin
        if(when_SuperResolutionPart3_l870) begin
          if(when_SuperResolutionPart3_l871) begin
            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_18[7:0];
          end else begin
            if(when_SuperResolutionPart3_l872) begin
              resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_20[7:0];
            end else begin
              resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_22[7:0];
            end
          end
        end else begin
          if(when_SuperResolutionPart3_l874) begin
            if(when_SuperResolutionPart3_l875) begin
              if(when_SuperResolutionPart3_l876) begin
                if(diffStage_controlPipe_payload_firstRow) begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_24[7:0];
                end else begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_26[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_28[7:0];
                  end
                end
              end else begin
                if(diffStage_controlPipe_payload_lastRow) begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_30[7:0];
                end else begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_32[7:0];
                end
              end
            end else begin
              if(when_SuperResolutionPart3_l884) begin
                if(when_SuperResolutionPart3_l885) begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_34[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_36[7:0];
                  end
                end else begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_38[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_40[7:0];
                  end
                end
              end else begin
                if(when_SuperResolutionPart3_l893) begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_42[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_44[7:0];
                  end
                end else begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_46[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_48[7:0];
                  end
                end
              end
            end
          end else begin
            if(when_SuperResolutionPart3_l902) begin
              if(when_SuperResolutionPart3_l903) begin
                if(diffStage_controlPipe_payload_firstRow) begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_50[7:0];
                end else begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_52[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_54[7:0];
                  end
                end
              end else begin
                if(diffStage_controlPipe_payload_lastRow) begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_56[7:0];
                end else begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_58[7:0];
                end
              end
            end else begin
              if(when_SuperResolutionPart3_l911) begin
                if(when_SuperResolutionPart3_l912) begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_60[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_62[7:0];
                  end
                end else begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_64[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_66[7:0];
                  end
                end
              end else begin
                if(when_SuperResolutionPart3_l920) begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_68[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_70[7:0];
                  end
                end else begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_72[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_74[7:0];
                  end
                end
              end
            end
          end
        end
      end else begin
        if(when_SuperResolutionPart3_l929) begin
          if(when_SuperResolutionPart3_l930) begin
            if(when_SuperResolutionPart3_l931) begin
              if(when_SuperResolutionPart3_l932) begin
                if(diffStage_controlPipe_payload_firstRow) begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_76[7:0];
                end else begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_78[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_80[7:0];
                  end
                end
              end else begin
                if(diffStage_controlPipe_payload_lastRow) begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_82[7:0];
                end else begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_84[7:0];
                end
              end
            end else begin
              if(when_SuperResolutionPart3_l940) begin
                if(when_SuperResolutionPart3_l941) begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_86[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_88[7:0];
                  end
                end else begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_90[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_92[7:0];
                  end
                end
              end else begin
                if(when_SuperResolutionPart3_l949) begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_94[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_96[7:0];
                  end
                end else begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_98[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_100[7:0];
                  end
                end
              end
            end
          end else begin
            if(when_SuperResolutionPart3_l958) begin
              if(when_SuperResolutionPart3_l959) begin
                if(diffStage_controlPipe_payload_firstRow) begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_102[7:0];
                end else begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_104[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_106[7:0];
                  end
                end
              end else begin
                if(diffStage_controlPipe_payload_lastRow) begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_108[7:0];
                end else begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_110[7:0];
                end
              end
            end else begin
              if(when_SuperResolutionPart3_l967) begin
                if(when_SuperResolutionPart3_l968) begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_112[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_114[7:0];
                  end
                end else begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_116[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_118[7:0];
                  end
                end
              end else begin
                if(when_SuperResolutionPart3_l976) begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_120[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_122[7:0];
                  end
                end else begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_124[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_126[7:0];
                  end
                end
              end
            end
          end
        end else begin
          if(when_SuperResolutionPart3_l985) begin
            if(when_SuperResolutionPart3_l986) begin
              if(when_SuperResolutionPart3_l987) begin
                resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_128[7:0];
              end else begin
                if(when_SuperResolutionPart3_l988) begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_130[7:0];
                end else begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_132[7:0];
                end
              end
            end else begin
              if(when_SuperResolutionPart3_l991) begin
                if(when_SuperResolutionPart3_l992) begin
                  if(diffStage_controlPipe_payload_firstRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_134[7:0];
                  end else begin
                    if(diffStage_controlPipe_payload_lastRow) begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_136[7:0];
                    end else begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_138[7:0];
                    end
                  end
                end else begin
                  if(diffStage_controlPipe_payload_lastRow) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_140[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_142[7:0];
                  end
                end
              end else begin
                if(when_SuperResolutionPart3_l1000) begin
                  if(when_SuperResolutionPart3_l1001) begin
                    if(diffStage_controlPipe_payload_lastRow) begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_144[7:0];
                    end else begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_146[7:0];
                    end
                  end else begin
                    if(diffStage_controlPipe_payload_lastRow) begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_148[7:0];
                    end else begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_150[7:0];
                    end
                  end
                end else begin
                  if(when_SuperResolutionPart3_l1009) begin
                    if(diffStage_controlPipe_payload_lastRow) begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_152[7:0];
                    end else begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_154[7:0];
                    end
                  end else begin
                    if(diffStage_controlPipe_payload_lastRow) begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_156[7:0];
                    end else begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_158[7:0];
                    end
                  end
                end
              end
            end
          end else begin
            if(when_SuperResolutionPart3_l1018) begin
              if(when_SuperResolutionPart3_l1019) begin
                if(when_SuperResolutionPart3_l1020) begin
                  resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_160[7:0];
                end else begin
                  if(when_SuperResolutionPart3_l1021) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_162[7:0];
                  end else begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_164[7:0];
                  end
                end
              end else begin
                if(when_SuperResolutionPart3_l1024) begin
                  if(when_SuperResolutionPart3_l1025) begin
                    if(diffStage_controlPipe_payload_firstRow) begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_166[7:0];
                    end else begin
                      if(diffStage_controlPipe_payload_lastRow) begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_168[7:0];
                      end else begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_170[7:0];
                      end
                    end
                  end else begin
                    if(diffStage_controlPipe_payload_lastRow) begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_172[7:0];
                    end else begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_174[7:0];
                    end
                  end
                end else begin
                  if(when_SuperResolutionPart3_l1033) begin
                    if(when_SuperResolutionPart3_l1034) begin
                      if(diffStage_controlPipe_payload_lastRow) begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_176[7:0];
                      end else begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_178[7:0];
                      end
                    end else begin
                      if(diffStage_controlPipe_payload_lastRow) begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_180[7:0];
                      end else begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_182[7:0];
                      end
                    end
                  end else begin
                    if(when_SuperResolutionPart3_l1042) begin
                      if(diffStage_controlPipe_payload_lastRow) begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_184[7:0];
                      end else begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_186[7:0];
                      end
                    end else begin
                      if(diffStage_controlPipe_payload_lastRow) begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_188[7:0];
                      end else begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_190[7:0];
                      end
                    end
                  end
                end
              end
            end else begin
              if(when_SuperResolutionPart3_l1051) begin
                if(when_SuperResolutionPart3_l1052) begin
                  if(when_SuperResolutionPart3_l1053) begin
                    if(diffStage_controlPipe_payload_firstRow) begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_192[7:0];
                    end else begin
                      if(diffStage_controlPipe_payload_lastRow) begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_194[7:0];
                      end else begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_196[7:0];
                      end
                    end
                  end else begin
                    if(diffStage_controlPipe_payload_lastRow) begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_198[7:0];
                    end else begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_200[7:0];
                    end
                  end
                end else begin
                  if(when_SuperResolutionPart3_l1061) begin
                    if(when_SuperResolutionPart3_l1062) begin
                      if(diffStage_controlPipe_payload_lastRow) begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_202[7:0];
                      end else begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_204[7:0];
                      end
                    end else begin
                      if(diffStage_controlPipe_payload_lastRow) begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_206[7:0];
                      end else begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_208[7:0];
                      end
                    end
                  end else begin
                    if(when_SuperResolutionPart3_l1070) begin
                      if(diffStage_controlPipe_payload_lastRow) begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_210[7:0];
                      end else begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_212[7:0];
                      end
                    end else begin
                      if(diffStage_controlPipe_payload_lastRow) begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_214[7:0];
                      end else begin
                        resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_216[7:0];
                      end
                    end
                  end
                end
              end else begin
                if(when_SuperResolutionPart3_l1078) begin
                  if(when_SuperResolutionPart3_l1079) begin
                    resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_218[7:0];
                  end else begin
                    if(when_SuperResolutionPart3_l1080) begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_220[7:0];
                    end else begin
                      resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_222[7:0];
                    end
                  end
                end else begin
                  if(when_SuperResolutionPart3_l1082) begin
                    if(when_SuperResolutionPart3_l1083) begin
                      if(when_SuperResolutionPart3_l1084) begin
                        if(diffStage_controlPipe_payload_firstRow) begin
                          resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_224[7:0];
                        end else begin
                          if(diffStage_controlPipe_payload_lastRow) begin
                            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_226[7:0];
                          end else begin
                            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_228[7:0];
                          end
                        end
                      end else begin
                        if(diffStage_controlPipe_payload_lastRow) begin
                          resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_230[7:0];
                        end else begin
                          resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_232[7:0];
                        end
                      end
                    end else begin
                      if(when_SuperResolutionPart3_l1092) begin
                        if(when_SuperResolutionPart3_l1093) begin
                          if(diffStage_controlPipe_payload_lastRow) begin
                            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_234[7:0];
                          end else begin
                            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_236[7:0];
                          end
                        end else begin
                          if(diffStage_controlPipe_payload_lastRow) begin
                            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_238[7:0];
                          end else begin
                            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_240[7:0];
                          end
                        end
                      end else begin
                        if(when_SuperResolutionPart3_l1101) begin
                          if(diffStage_controlPipe_payload_lastRow) begin
                            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_242[7:0];
                          end else begin
                            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_244[7:0];
                          end
                        end else begin
                          if(diffStage_controlPipe_payload_lastRow) begin
                            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_246[7:0];
                          end else begin
                            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_248[7:0];
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
  end

  assign when_SuperResolutionPart3_l840 = ((diffStage_controlPipe_payload_currentPosition == 2'b00) && diffStage_mainOneValidStream_payload);
  assign when_SuperResolutionPart3_l846 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l847 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l850 = (minDiff < diffStage_controlPipe_payload_verticalDiff);
  assign when_SuperResolutionPart3_l854 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l855 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l860 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l861 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l851 = (diffStage_controlPipe_payload_verticalDiff == minDiff);
  assign when_SuperResolutionPart3_l841 = ((diffStage_controlPipe_payload_currentPosition == 2'b01) && diffStage_mainTwoValidStream_payload);
  assign when_SuperResolutionPart3_l842 = ((diffStage_controlPipe_payload_currentPosition == 2'b10) && diffStage_mainThreeValidStream_payload);
  assign when_SuperResolutionPart3_l869 = ((diffStage_controlPipe_payload_horizontalDirectionValid && diffStage_controlPipe_payload_mainDirectionValid) && diffStage_controlPipe_payload_counterDirectionValid);
  assign when_SuperResolutionPart3_l870 = ((diffStage_controlPipe_payload_horizontalDiff <= diffStage_controlPipe_payload_mainDiff) && (diffStage_controlPipe_payload_horizontalDiff <= diffStage_controlPipe_payload_counterDiff));
  assign when_SuperResolutionPart3_l871 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l872 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l875 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l876 = (diffStage_controlPipe_payload_nextPosition == 2'b01);
  assign when_SuperResolutionPart3_l885 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l893 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l884 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l902 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l903 = (diffStage_controlPipe_payload_nextPosition == 2'b01);
  assign when_SuperResolutionPart3_l912 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l920 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l911 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l874 = ((diffStage_controlPipe_payload_mainDiff < diffStage_controlPipe_payload_horizontalDiff) && (diffStage_controlPipe_payload_mainDiff <= diffStage_controlPipe_payload_counterDiff));
  assign when_SuperResolutionPart3_l930 = (diffStage_controlPipe_payload_mainDiff <= diffStage_controlPipe_payload_counterDiff);
  assign when_SuperResolutionPart3_l931 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l932 = (diffStage_controlPipe_payload_nextPosition == 2'b01);
  assign when_SuperResolutionPart3_l941 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l949 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l940 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l958 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l959 = (diffStage_controlPipe_payload_nextPosition == 2'b01);
  assign when_SuperResolutionPart3_l968 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l976 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l967 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l986 = (diffStage_controlPipe_payload_horizontalDiff <= diffStage_controlPipe_payload_counterDiff);
  assign when_SuperResolutionPart3_l987 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l988 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l991 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l992 = (diffStage_controlPipe_payload_nextPosition == 2'b01);
  assign when_SuperResolutionPart3_l1001 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l1009 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l1000 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l1019 = (diffStage_controlPipe_payload_horizontalDiff <= diffStage_controlPipe_payload_mainDiff);
  assign when_SuperResolutionPart3_l1020 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l1021 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l1024 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l1025 = (diffStage_controlPipe_payload_nextPosition == 2'b01);
  assign when_SuperResolutionPart3_l1034 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l1042 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l1033 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l1052 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l1053 = (diffStage_controlPipe_payload_nextPosition == 2'b01);
  assign when_SuperResolutionPart3_l1062 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l1070 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l1061 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l1079 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l1080 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l1083 = (diffStage_controlPipe_payload_currentPosition == 2'b00);
  assign when_SuperResolutionPart3_l1084 = (diffStage_controlPipe_payload_nextPosition == 2'b01);
  assign when_SuperResolutionPart3_l1093 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l1101 = (diffStage_controlPipe_payload_nextPosition == 2'b00);
  assign when_SuperResolutionPart3_l1092 = (diffStage_controlPipe_payload_currentPosition == 2'b01);
  assign when_SuperResolutionPart3_l929 = (((! diffStage_controlPipe_payload_horizontalDirectionValid) && diffStage_controlPipe_payload_mainDirectionValid) && diffStage_controlPipe_payload_counterDirectionValid);
  assign when_SuperResolutionPart3_l985 = ((diffStage_controlPipe_payload_horizontalDirectionValid && (! diffStage_controlPipe_payload_mainDirectionValid)) && diffStage_controlPipe_payload_counterDirectionValid);
  assign when_SuperResolutionPart3_l1018 = ((diffStage_controlPipe_payload_horizontalDirectionValid && diffStage_controlPipe_payload_mainDirectionValid) && (! diffStage_controlPipe_payload_counterDirectionValid));
  assign when_SuperResolutionPart3_l1051 = (((! diffStage_controlPipe_payload_horizontalDirectionValid) && (! diffStage_controlPipe_payload_mainDirectionValid)) && diffStage_controlPipe_payload_counterDirectionValid);
  assign when_SuperResolutionPart3_l1078 = ((diffStage_controlPipe_payload_horizontalDirectionValid && (! diffStage_controlPipe_payload_mainDirectionValid)) && (! diffStage_controlPipe_payload_counterDirectionValid));
  assign when_SuperResolutionPart3_l1082 = (((! diffStage_controlPipe_payload_horizontalDirectionValid) && diffStage_controlPipe_payload_mainDirectionValid) && (! diffStage_controlPipe_payload_counterDirectionValid));
  assign resultStage_pixelStream_ready = (! resultStage_pixelStream_rValid);
  assign resultStage_pixelStream_s2mPipe_valid = (resultStage_pixelStream_valid || resultStage_pixelStream_rValid);
  assign resultStage_pixelStream_s2mPipe_payload = (resultStage_pixelStream_rValid ? resultStage_pixelStream_rData : resultStage_pixelStream_payload);
  always @(*) begin
    resultStage_pixelStream_s2mPipe_ready = resultStage_resultStream_ready;
    if(when_Stream_l368_67) begin
      resultStage_pixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_67 = (! resultStage_resultStream_valid);
  assign resultStage_resultStream_valid = resultStage_pixelStream_s2mPipe_rValid;
  assign resultStage_resultStream_payload = resultStage_pixelStream_s2mPipe_rData;
  assign when_SuperResolutionPart3_l1115 = (! resultStage_controlPipeBeforePipe_payload_finalResult);
  assign diffStage_controlPipe_fire = (diffStage_controlPipe_valid && diffStage_controlPipe_ready);
  assign CICC1851_resultStage_mainOnePixelStream_ready_2 = (CICC1851_resultStage_mainOnePixelStream_ready && CICC1851_resultStage_mainOnePixelStream_ready_1);
  assign CICC1851_resultStage_mainOnePixelStream_ready = (((((((((((((resultStage_resultStream_valid && resultStage_mainOnePixelStream_valid) && resultStage_counterOnePixelStream_valid) && resultStage_mainTwoPixelStream_valid) && resultStage_counterTwoPixelStream_valid) && resultStage_mainThreePixelStream_valid) && resultStage_counterThreePixelStream_valid) && resultStage_mainOneValidStream_valid) && resultStage_counterOneValidStream_valid) && resultStage_mainTwoValidStream_valid) && resultStage_counterTwoValidStream_valid) && resultStage_mainThreeValidStream_valid) && resultStage_counterThreeValidStream_valid) && resultStage_controlPipe_valid);
  assign resultStage_resultStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_mainOnePixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_counterOnePixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_mainTwoPixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_counterTwoPixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_mainThreePixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_counterThreePixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_mainOneValidStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_counterOneValidStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_mainTwoValidStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_counterTwoValidStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_mainThreeValidStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_counterThreeValidStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_controlPipe_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign when_Stream_l438 = ((! resultStage_controlPipe_payload_pipeValid) || (! resultStage_controlPipe_payload_finalResult));
  always @(*) begin
    resultsJoin_valid = CICC1851_resultStage_mainOnePixelStream_ready;
    if(when_Stream_l438) begin
      resultsJoin_valid = 1'b0;
    end
  end

  always @(*) begin
    CICC1851_resultStage_mainOnePixelStream_ready_1 = resultsJoin_ready;
    if(when_Stream_l438) begin
      CICC1851_resultStage_mainOnePixelStream_ready_1 = 1'b1;
    end
  end

  assign pixelsStream_valid = resultsJoin_valid;
  assign resultsJoin_ready = pixelsStream_ready;
  assign pixelsStream_payload_pixel = resultStage_resultStream_payload;
  assign pixelsStream_payload_frameStart = resultStage_controlPipe_payload_frameStart;
  assign pixelsStream_payload_rowEnd = resultStage_controlPipe_payload_rowEnd;
  assign pixelsStream_ready = (! pixelsStream_rValid);
  assign pixelsStream_s2mPipe_valid = (pixelsStream_valid || pixelsStream_rValid);
  assign pixelsStream_s2mPipe_payload_pixel = (pixelsStream_rValid ? pixelsStream_rData_pixel : pixelsStream_payload_pixel);
  assign pixelsStream_s2mPipe_payload_frameStart = (pixelsStream_rValid ? pixelsStream_rData_frameStart : pixelsStream_payload_frameStart);
  assign pixelsStream_s2mPipe_payload_rowEnd = (pixelsStream_rValid ? pixelsStream_rData_rowEnd : pixelsStream_payload_rowEnd);
  always @(*) begin
    pixelsStream_s2mPipe_ready = pixelsStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_68) begin
      pixelsStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_68 = (! pixelsStream_s2mPipe_m2sPipe_valid);
  assign pixelsStream_s2mPipe_m2sPipe_valid = pixelsStream_s2mPipe_rValid;
  assign pixelsStream_s2mPipe_m2sPipe_payload_pixel = pixelsStream_s2mPipe_rData_pixel;
  assign pixelsStream_s2mPipe_m2sPipe_payload_frameStart = pixelsStream_s2mPipe_rData_frameStart;
  assign pixelsStream_s2mPipe_m2sPipe_payload_rowEnd = pixelsStream_s2mPipe_rData_rowEnd;
  assign pixelsStream_s2mPipe_m2sPipe_ready = pixelsOut_ready;
  assign controlStateMachine_wantExit = 1'b0;
  always @(*) begin
    controlStateMachine_wantStart = 1'b0;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_2_HOLD : begin
      end
      controlStateMachine_enumDef_2_PASS : begin
      end
      controlStateMachine_enumDef_2_EXTRA : begin
      end
      default : begin
        controlStateMachine_wantStart = 1'b1;
      end
    endcase
  end

  assign controlStateMachine_wantKill = 1'b0;
  always @(*) begin
    controlStateMachine_stateNext = controlStateMachine_stateReg;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_2_HOLD : begin
        if(passPixels_fire_13) begin
          if(when_SuperResolutionPart3_l1158) begin
            controlStateMachine_stateNext = controlStateMachine_enumDef_2_PASS;
          end
        end
      end
      controlStateMachine_enumDef_2_PASS : begin
        if(controlStream_fire) begin
          controlStateMachine_stateNext = controlStateMachine_enumDef_2_EXTRA;
        end
      end
      controlStateMachine_enumDef_2_EXTRA : begin
        if(controlStream_fire_1) begin
          if(writeDone) begin
            if(when_SuperResolutionPart3_l1199) begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_2_HOLD;
            end else begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_2_PASS;
            end
          end else begin
            if(outReachRowEnd) begin
              if(when_SuperResolutionPart3_l1202) begin
                controlStateMachine_stateNext = controlStateMachine_enumDef_2_PASS;
              end else begin
                controlStateMachine_stateNext = controlStateMachine_enumDef_2_HOLD;
              end
            end else begin
              if(when_SuperResolutionPart3_l1205) begin
                controlStateMachine_stateNext = controlStateMachine_enumDef_2_PASS;
              end else begin
                controlStateMachine_stateNext = controlStateMachine_enumDef_2_HOLD;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
    if(controlStateMachine_wantStart) begin
      controlStateMachine_stateNext = controlStateMachine_enumDef_2_HOLD;
    end
    if(controlStateMachine_wantKill) begin
      controlStateMachine_stateNext = controlStateMachine_enumDef_2_BOOT;
    end
  end

  assign passPixels_fire_13 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart3_l1158 = ((outRowCount_value < bufferRowCount_value) && (outPixelAddr_value < bufferWAddr_value));
  assign controlStream_fire = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart3_l1168 = (outPixelAddr_value == 12'h0);
  assign when_SuperResolutionPart3_l1188 = (outRowCount_value == 12'h0);
  assign controlStream_fire_1 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart3_l1199 = (outReachFinalRow && outReachRowEnd);
  assign passPixels_fire_14 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart3_l1202 = (((bufferRowCount_value == CICC1851_when_SuperResolutionPart3_l1202) || (12'h001 < bufferWAddr_value)) || ((bufferWAddr_value == 12'h001) && passPixels_fire_14));
  assign passPixels_fire_15 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart3_l1205 = (((CICC1851_when_SuperResolutionPart3_l1205 < bufferRowCount_value) || ((bufferWAddr_value == CICC1851_when_SuperResolutionPart3_l1205_1) && passPixels_fire_15)) || (CICC1851_when_SuperResolutionPart3_l1205_2 < bufferWAddr_value));
  assign when_SuperResolutionPart3_l1217 = (outRowCount_value == 12'h0);
  assign controlStream_fire_2 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart3_l1220 = (frameStart && controlStream_fire_2);
  assign controlStream_fire_3 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart3_l1223 = (controlStream_fire_3 && (CICC1851_when_SuperResolutionPart3_l1223 == CICC1851_when_SuperResolutionPart3_l1223_1));
  assign controlStream_fire_4 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart3_l1224 = ((outReachRowEnd && (CICC1851_when_SuperResolutionPart3_l1224 == CICC1851_when_SuperResolutionPart3_l1224_1)) && controlStream_fire_4);
  assign controlStream_fire_5 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart3_l1226 = (controlStream_fire_5 && outReachRowEnd);
  assign controlStream_fire_6 = (controlStream_valid && controlStream_ready);
  assign controlStream_fire_7 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart3_l1247 = (controlStream_payload_rowEnd && controlStream_fire_7);
  assign when_SuperResolutionPart3_l1248 = (outRowCount_value != 12'h0);
  assign when_SuperResolutionPart3_l1250 = (currentRowBuffer == 2'b10);
  assign when_SuperResolutionPart3_l1252 = (nextRowBuffer == 2'b10);
  always @(posedge clk or negedge resetn) begin
    if(!resetn) begin
      inpThreeDone <= 1'b0;
      readDone <= 1'b0;
      startRead <= 1'b0;
      frameStart <= 1'b0;
      inpThreshold <= 8'h80;
      bmpWidth <= 10'h3c0;
      bmpHeight <= 10'h21c;
      holdBuffer <= 1'b0;
      writeDone <= 1'b0;
      bufferRowCount_value <= 12'h0;
      bufferEnable <= 1'b0;
      bufferSwitch <= 2'b00;
      nextRowBuffer <= 2'b01;
      currentRowBuffer <= 2'b00;
      bufferReuse <= 1'b0;
      bufferWAddr_value <= 12'h0;
      outPixelAddr_value <= 12'h0;
      outRowCount_value <= 12'h0;
      alreadySendRow_value <= 12'h0;
      alreadySendCountInRow_value <= 12'h0;
      alreadyReachRowEnd <= 1'b0;
      alreadyReachFinalRow <= 1'b0;
      outReachRowEnd <= 1'b0;
      outReachFinalRow <= 1'b0;
      bufferReachRowEnd <= 1'b0;
      bufferReachFinalRow <= 1'b0;
      minDiff <= 8'h0;
      candidatePixel <= 8'h0;
      isHorizontalDirection <= 1'b0;
      inValidMinDiff <= 1'b0;
      pixelsIn_rValid <= 1'b0;
      pixelsIn_s2mPipe_rValid <= 1'b0;
      mainPixelAddrOneStream_rValid <= 1'b0;
      mainPixelAddrOneStream_s2mPipe_rValid <= 1'b0;
      CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_mainOnePixelStream_valid <= 1'b0;
      counterPixelAddrOneStream_rValid <= 1'b0;
      counterPixelAddrOneStream_s2mPipe_rValid <= 1'b0;
      CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_counterOnePixelStream_valid <= 1'b0;
      mainPixelAddrTwoStream_rValid <= 1'b0;
      mainPixelAddrTwoStream_s2mPipe_rValid <= 1'b0;
      CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_mainTwoPixelStream_valid <= 1'b0;
      counterPixelAddrTwoStream_rValid <= 1'b0;
      counterPixelAddrTwoStream_s2mPipe_rValid <= 1'b0;
      CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_counterTwoPixelStream_valid <= 1'b0;
      mainPixelAddrThreeStream_rValid <= 1'b0;
      mainPixelAddrThreeStream_s2mPipe_rValid <= 1'b0;
      CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_mainThreePixelStream_valid <= 1'b0;
      counterPixelAddrThreeStream_rValid <= 1'b0;
      counterPixelAddrThreeStream_s2mPipe_rValid <= 1'b0;
      CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_counterThreePixelStream_valid <= 1'b0;
      mainValidAddrOneStream_rValid <= 1'b0;
      mainValidAddrOneStream_s2mPipe_rValid <= 1'b0;
      CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_mainOneValidStream_valid <= 1'b0;
      counterValidAddrOneStream_rValid <= 1'b0;
      counterValidAddrOneStream_s2mPipe_rValid <= 1'b0;
      CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_counterOneValidStream_valid <= 1'b0;
      mainValidAddrTwoStream_rValid <= 1'b0;
      mainValidAddrTwoStream_s2mPipe_rValid <= 1'b0;
      CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_mainTwoValidStream_valid <= 1'b0;
      counterValidAddrTwoStream_rValid <= 1'b0;
      counterValidAddrTwoStream_s2mPipe_rValid <= 1'b0;
      CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_counterTwoValidStream_valid <= 1'b0;
      mainValidAddrThreeStream_rValid <= 1'b0;
      mainValidAddrThreeStream_s2mPipe_rValid <= 1'b0;
      CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_mainThreeValidStream_valid <= 1'b0;
      counterValidAddrThreeStream_rValid <= 1'b0;
      counterValidAddrThreeStream_s2mPipe_rValid <= 1'b0;
      CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_counterThreeValidStream_valid <= 1'b0;
      controlStream_rValid <= 1'b0;
      controlStream_s2mPipe_rValid <= 1'b0;
      controlStream_s2mPipe_m2sPipe_rValid <= 1'b0;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rValid <= 1'b0;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rValid <= 1'b0;
      readStage_mainOnePixelStream_rValid <= 1'b0;
      readStage_mainOnePixelStream_s2mPipe_rValid <= 1'b0;
      readStage_counterOnePixelStream_rValid <= 1'b0;
      readStage_counterOnePixelStream_s2mPipe_rValid <= 1'b0;
      readStage_mainTwoPixelStream_rValid <= 1'b0;
      readStage_mainTwoPixelStream_s2mPipe_rValid <= 1'b0;
      readStage_counterTwoPixelStream_rValid <= 1'b0;
      readStage_counterTwoPixelStream_s2mPipe_rValid <= 1'b0;
      readStage_mainThreePixelStream_rValid <= 1'b0;
      readStage_mainThreePixelStream_s2mPipe_rValid <= 1'b0;
      readStage_counterThreePixelStream_rValid <= 1'b0;
      readStage_counterThreePixelStream_s2mPipe_rValid <= 1'b0;
      readStage_mainOneValidStream_rValid <= 1'b0;
      readStage_mainOneValidStream_s2mPipe_rValid <= 1'b0;
      readStage_counterOneValidStream_rValid <= 1'b0;
      readStage_counterOneValidStream_s2mPipe_rValid <= 1'b0;
      readStage_mainTwoValidStream_rValid <= 1'b0;
      readStage_mainTwoValidStream_s2mPipe_rValid <= 1'b0;
      readStage_counterTwoValidStream_rValid <= 1'b0;
      readStage_counterTwoValidStream_s2mPipe_rValid <= 1'b0;
      readStage_mainThreeValidStream_rValid <= 1'b0;
      readStage_mainThreeValidStream_s2mPipe_rValid <= 1'b0;
      readStage_counterThreeValidStream_rValid <= 1'b0;
      readStage_counterThreeValidStream_s2mPipe_rValid <= 1'b0;
      readStage_controlPipe_translated_rValid <= 1'b0;
      readStage_controlPipe_translated_s2mPipe_rValid <= 1'b0;
      compareStage_mainOnePixelStream_rValid <= 1'b0;
      compareStage_mainOnePixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_counterOnePixelStream_rValid <= 1'b0;
      compareStage_counterOnePixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_mainTwoPixelStream_rValid <= 1'b0;
      compareStage_mainTwoPixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_counterTwoPixelStream_rValid <= 1'b0;
      compareStage_counterTwoPixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_mainThreePixelStream_rValid <= 1'b0;
      compareStage_mainThreePixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_counterThreePixelStream_rValid <= 1'b0;
      compareStage_counterThreePixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_mainOneValidStream_rValid <= 1'b0;
      compareStage_mainOneValidStream_s2mPipe_rValid <= 1'b0;
      compareStage_counterOneValidStream_rValid <= 1'b0;
      compareStage_counterOneValidStream_s2mPipe_rValid <= 1'b0;
      compareStage_mainTwoValidStream_rValid <= 1'b0;
      compareStage_mainTwoValidStream_s2mPipe_rValid <= 1'b0;
      compareStage_counterTwoValidStream_rValid <= 1'b0;
      compareStage_counterTwoValidStream_s2mPipe_rValid <= 1'b0;
      compareStage_mainThreeValidStream_rValid <= 1'b0;
      compareStage_mainThreeValidStream_s2mPipe_rValid <= 1'b0;
      compareStage_counterThreeValidStream_rValid <= 1'b0;
      compareStage_counterThreeValidStream_s2mPipe_rValid <= 1'b0;
      compareStage_controlPipe_translated_rValid <= 1'b0;
      compareStage_controlPipe_translated_s2mPipe_rValid <= 1'b0;
      diffStage_mainOnePixelStream_rValid <= 1'b0;
      diffStage_mainOnePixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_counterOnePixelStream_rValid <= 1'b0;
      diffStage_counterOnePixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_mainTwoPixelStream_rValid <= 1'b0;
      diffStage_mainTwoPixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_counterTwoPixelStream_rValid <= 1'b0;
      diffStage_counterTwoPixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_mainThreePixelStream_rValid <= 1'b0;
      diffStage_mainThreePixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_counterThreePixelStream_rValid <= 1'b0;
      diffStage_counterThreePixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_mainOneValidStream_rValid <= 1'b0;
      diffStage_mainOneValidStream_s2mPipe_rValid <= 1'b0;
      diffStage_counterOneValidStream_rValid <= 1'b0;
      diffStage_counterOneValidStream_s2mPipe_rValid <= 1'b0;
      diffStage_mainTwoValidStream_rValid <= 1'b0;
      diffStage_mainTwoValidStream_s2mPipe_rValid <= 1'b0;
      diffStage_counterTwoValidStream_rValid <= 1'b0;
      diffStage_counterTwoValidStream_s2mPipe_rValid <= 1'b0;
      diffStage_mainThreeValidStream_rValid <= 1'b0;
      diffStage_mainThreeValidStream_s2mPipe_rValid <= 1'b0;
      diffStage_counterThreeValidStream_rValid <= 1'b0;
      diffStage_counterThreeValidStream_s2mPipe_rValid <= 1'b0;
      resultStage_controlPipeBeforePipe_rValid <= 1'b0;
      resultStage_controlPipeBeforePipe_s2mPipe_rValid <= 1'b0;
      resultStage_pixelStream_rValid <= 1'b0;
      resultStage_pixelStream_s2mPipe_rValid <= 1'b0;
      pixelsStream_rValid <= 1'b0;
      pixelsStream_s2mPipe_rValid <= 1'b0;
      controlStateMachine_stateReg <= controlStateMachine_enumDef_2_BOOT;
    end else begin
      if(when_SuperResolutionPart3_l72) begin
        inpThreeDone <= 1'b0;
      end
      if(when_SuperResolutionPart3_l75) begin
        readDone <= 1'b0;
      end
      if(when_SuperResolutionPart3_l78) begin
        startRead <= 1'b1;
      end
      if(when_SuperResolutionPart3_l78_1) begin
        startRead <= 1'b0;
      end
      inpThreshold <= thresholdIn;
      bmpWidth <= widthIn;
      bmpHeight <= heightIn;
      if(when_SuperResolutionPart3_l93) begin
        holdBuffer <= 1'b0;
      end
      if(when_SuperResolutionPart3_l96) begin
        writeDone <= 1'b0;
      end
      bufferRowCount_value <= bufferRowCount_valueNext;
      if(when_SuperResolutionPart3_l102) begin
        bufferEnable <= 1'b1;
      end
      if(when_SuperResolutionPart3_l102_1) begin
        bufferEnable <= 1'b0;
      end
      if(inpThreeDone) begin
        bufferReuse <= 1'b0;
      end
      bufferWAddr_value <= bufferWAddr_valueNext;
      outPixelAddr_value <= outPixelAddr_valueNext;
      outRowCount_value <= outRowCount_valueNext;
      alreadySendRow_value <= alreadySendRow_valueNext;
      alreadySendCountInRow_value <= alreadySendCountInRow_valueNext;
      if(when_SuperResolutionPart3_l154) begin
        bufferSwitch <= 2'b00;
        nextRowBuffer <= {1'd0, CICC1851_nextRowBuffer};
        currentRowBuffer <= 2'b00;
        minDiff <= 8'h0;
        candidatePixel <= 8'h0;
        isHorizontalDirection <= 1'b0;
      end
      if(pixelsIn_valid) begin
        pixelsIn_rValid <= 1'b1;
      end
      if(pixelsIn_s2mPipe_ready) begin
        pixelsIn_rValid <= 1'b0;
      end
      if(pixelsIn_s2mPipe_ready) begin
        pixelsIn_s2mPipe_rValid <= pixelsIn_s2mPipe_valid;
      end
      if(when_SuperResolutionPart3_l226) begin
        bufferReachRowEnd <= 1'b1;
      end
      if(when_SuperResolutionPart3_l227) begin
        bufferReachFinalRow <= 1'b1;
      end
      if(when_SuperResolutionPart3_l230) begin
        if(bufferReachFinalRow) begin
          bufferReuse <= 1'b1;
          bufferReachRowEnd <= 1'b0;
          bufferReachFinalRow <= 1'b0;
        end else begin
          bufferReachRowEnd <= 1'b0;
        end
      end
      if(when_SuperResolutionPart3_l243) begin
        if(when_SuperResolutionPart3_l244) begin
          bufferSwitch <= 2'b00;
        end else begin
          bufferSwitch <= (bufferSwitch + 2'b01);
        end
      end
      if(when_SuperResolutionPart3_l251) begin
        holdBuffer <= 1'b1;
        bufferEnable <= 1'b0;
        if(when_SuperResolutionPart3_l255) begin
          writeDone <= 1'b1;
          bufferEnable <= 1'b0;
        end
      end
      if(when_SuperResolutionPart3_l262) begin
        frameStart <= 1'b1;
      end
      if(inpThreeDone) begin
        inpThreeDone <= 1'b0;
      end
      if(when_SuperResolutionPart3_l270) begin
        alreadyReachRowEnd <= 1'b1;
      end
      if(when_SuperResolutionPart3_l271) begin
        alreadyReachFinalRow <= 1'b1;
      end
      if(pixelsOut_fire_2) begin
        if(alreadyReachRowEnd) begin
          alreadyReachRowEnd <= 1'b0;
          if(alreadyReachFinalRow) begin
            alreadyReachFinalRow <= 1'b0;
          end
        end
      end
      if(when_SuperResolutionPart3_l282) begin
        inpThreeDone <= 1'b1;
      end
      if(mainPixelAddrOneStream_valid) begin
        mainPixelAddrOneStream_rValid <= 1'b1;
      end
      if(mainPixelAddrOneStream_s2mPipe_ready) begin
        mainPixelAddrOneStream_rValid <= 1'b0;
      end
      if(mainPixelAddrOneStream_s2mPipe_ready) begin
        mainPixelAddrOneStream_s2mPipe_rValid <= mainPixelAddrOneStream_s2mPipe_valid;
      end
      if(CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(mainPixelAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_2 <= mainPixelAddrOneStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_1) begin
        CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_1) begin
        CICC1851_readStage_mainOnePixelStream_valid <= (CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready || CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_3);
      end
      if(counterPixelAddrOneStream_valid) begin
        counterPixelAddrOneStream_rValid <= 1'b1;
      end
      if(counterPixelAddrOneStream_s2mPipe_ready) begin
        counterPixelAddrOneStream_rValid <= 1'b0;
      end
      if(counterPixelAddrOneStream_s2mPipe_ready) begin
        counterPixelAddrOneStream_s2mPipe_rValid <= counterPixelAddrOneStream_s2mPipe_valid;
      end
      if(CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(counterPixelAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_2 <= counterPixelAddrOneStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_2) begin
        CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_2) begin
        CICC1851_readStage_counterOnePixelStream_valid <= (CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready || CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_3);
      end
      if(mainPixelAddrTwoStream_valid) begin
        mainPixelAddrTwoStream_rValid <= 1'b1;
      end
      if(mainPixelAddrTwoStream_s2mPipe_ready) begin
        mainPixelAddrTwoStream_rValid <= 1'b0;
      end
      if(mainPixelAddrTwoStream_s2mPipe_ready) begin
        mainPixelAddrTwoStream_s2mPipe_rValid <= mainPixelAddrTwoStream_s2mPipe_valid;
      end
      if(CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= mainPixelAddrTwoStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_3) begin
        CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_3) begin
        CICC1851_readStage_mainTwoPixelStream_valid <= (CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready || CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_3);
      end
      if(counterPixelAddrTwoStream_valid) begin
        counterPixelAddrTwoStream_rValid <= 1'b1;
      end
      if(counterPixelAddrTwoStream_s2mPipe_ready) begin
        counterPixelAddrTwoStream_rValid <= 1'b0;
      end
      if(counterPixelAddrTwoStream_s2mPipe_ready) begin
        counterPixelAddrTwoStream_s2mPipe_rValid <= counterPixelAddrTwoStream_s2mPipe_valid;
      end
      if(CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= counterPixelAddrTwoStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_4) begin
        CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_4) begin
        CICC1851_readStage_counterTwoPixelStream_valid <= (CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready || CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_3);
      end
      if(mainPixelAddrThreeStream_valid) begin
        mainPixelAddrThreeStream_rValid <= 1'b1;
      end
      if(mainPixelAddrThreeStream_s2mPipe_ready) begin
        mainPixelAddrThreeStream_rValid <= 1'b0;
      end
      if(mainPixelAddrThreeStream_s2mPipe_ready) begin
        mainPixelAddrThreeStream_s2mPipe_rValid <= mainPixelAddrThreeStream_s2mPipe_valid;
      end
      if(CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_2 <= mainPixelAddrThreeStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_5) begin
        CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_5) begin
        CICC1851_readStage_mainThreePixelStream_valid <= (CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready || CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_3);
      end
      if(counterPixelAddrThreeStream_valid) begin
        counterPixelAddrThreeStream_rValid <= 1'b1;
      end
      if(counterPixelAddrThreeStream_s2mPipe_ready) begin
        counterPixelAddrThreeStream_rValid <= 1'b0;
      end
      if(counterPixelAddrThreeStream_s2mPipe_ready) begin
        counterPixelAddrThreeStream_s2mPipe_rValid <= counterPixelAddrThreeStream_s2mPipe_valid;
      end
      if(CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_2 <= counterPixelAddrThreeStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_6) begin
        CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_6) begin
        CICC1851_readStage_counterThreePixelStream_valid <= (CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready || CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_3);
      end
      if(mainValidAddrOneStream_valid) begin
        mainValidAddrOneStream_rValid <= 1'b1;
      end
      if(mainValidAddrOneStream_s2mPipe_ready) begin
        mainValidAddrOneStream_rValid <= 1'b0;
      end
      if(mainValidAddrOneStream_s2mPipe_ready) begin
        mainValidAddrOneStream_s2mPipe_rValid <= mainValidAddrOneStream_s2mPipe_valid;
      end
      if(CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(mainValidAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_2 <= mainValidAddrOneStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_7) begin
        CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_7) begin
        CICC1851_readStage_mainOneValidStream_valid <= (CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready || CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_3);
      end
      if(counterValidAddrOneStream_valid) begin
        counterValidAddrOneStream_rValid <= 1'b1;
      end
      if(counterValidAddrOneStream_s2mPipe_ready) begin
        counterValidAddrOneStream_rValid <= 1'b0;
      end
      if(counterValidAddrOneStream_s2mPipe_ready) begin
        counterValidAddrOneStream_s2mPipe_rValid <= counterValidAddrOneStream_s2mPipe_valid;
      end
      if(CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(counterValidAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_2 <= counterValidAddrOneStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_8) begin
        CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_8) begin
        CICC1851_readStage_counterOneValidStream_valid <= (CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready || CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_3);
      end
      if(mainValidAddrTwoStream_valid) begin
        mainValidAddrTwoStream_rValid <= 1'b1;
      end
      if(mainValidAddrTwoStream_s2mPipe_ready) begin
        mainValidAddrTwoStream_rValid <= 1'b0;
      end
      if(mainValidAddrTwoStream_s2mPipe_ready) begin
        mainValidAddrTwoStream_s2mPipe_rValid <= mainValidAddrTwoStream_s2mPipe_valid;
      end
      if(CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(mainValidAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= mainValidAddrTwoStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_9) begin
        CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_9) begin
        CICC1851_readStage_mainTwoValidStream_valid <= (CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready || CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_3);
      end
      if(counterValidAddrTwoStream_valid) begin
        counterValidAddrTwoStream_rValid <= 1'b1;
      end
      if(counterValidAddrTwoStream_s2mPipe_ready) begin
        counterValidAddrTwoStream_rValid <= 1'b0;
      end
      if(counterValidAddrTwoStream_s2mPipe_ready) begin
        counterValidAddrTwoStream_s2mPipe_rValid <= counterValidAddrTwoStream_s2mPipe_valid;
      end
      if(CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(counterValidAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= counterValidAddrTwoStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_10) begin
        CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_10) begin
        CICC1851_readStage_counterTwoValidStream_valid <= (CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready || CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_3);
      end
      if(mainValidAddrThreeStream_valid) begin
        mainValidAddrThreeStream_rValid <= 1'b1;
      end
      if(mainValidAddrThreeStream_s2mPipe_ready) begin
        mainValidAddrThreeStream_rValid <= 1'b0;
      end
      if(mainValidAddrThreeStream_s2mPipe_ready) begin
        mainValidAddrThreeStream_s2mPipe_rValid <= mainValidAddrThreeStream_s2mPipe_valid;
      end
      if(CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(mainValidAddrThreeStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_2 <= mainValidAddrThreeStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_11) begin
        CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_11) begin
        CICC1851_readStage_mainThreeValidStream_valid <= (CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready || CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_3);
      end
      if(counterValidAddrThreeStream_valid) begin
        counterValidAddrThreeStream_rValid <= 1'b1;
      end
      if(counterValidAddrThreeStream_s2mPipe_ready) begin
        counterValidAddrThreeStream_rValid <= 1'b0;
      end
      if(counterValidAddrThreeStream_s2mPipe_ready) begin
        counterValidAddrThreeStream_s2mPipe_rValid <= counterValidAddrThreeStream_s2mPipe_valid;
      end
      if(CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(counterValidAddrThreeStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_2 <= counterValidAddrThreeStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_12) begin
        CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_12) begin
        CICC1851_readStage_counterThreeValidStream_valid <= (CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready || CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_3);
      end
      if(controlStream_valid) begin
        controlStream_rValid <= 1'b1;
      end
      if(controlStream_s2mPipe_ready) begin
        controlStream_rValid <= 1'b0;
      end
      if(controlStream_s2mPipe_ready) begin
        controlStream_s2mPipe_rValid <= controlStream_s2mPipe_valid;
      end
      if(controlStream_s2mPipe_m2sPipe_ready) begin
        controlStream_s2mPipe_m2sPipe_rValid <= controlStream_s2mPipe_m2sPipe_valid;
      end
      if(controlStream_s2mPipe_m2sPipe_m2sPipe_valid) begin
        controlStream_s2mPipe_m2sPipe_m2sPipe_rValid <= 1'b1;
      end
      if(controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready) begin
        controlStream_s2mPipe_m2sPipe_m2sPipe_rValid <= 1'b0;
      end
      if(controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready) begin
        controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_valid;
      end
      if(readStage_mainOnePixelStream_valid) begin
        readStage_mainOnePixelStream_rValid <= 1'b1;
      end
      if(readStage_mainOnePixelStream_s2mPipe_ready) begin
        readStage_mainOnePixelStream_rValid <= 1'b0;
      end
      if(readStage_mainOnePixelStream_s2mPipe_ready) begin
        readStage_mainOnePixelStream_s2mPipe_rValid <= readStage_mainOnePixelStream_s2mPipe_valid;
      end
      if(readStage_counterOnePixelStream_valid) begin
        readStage_counterOnePixelStream_rValid <= 1'b1;
      end
      if(readStage_counterOnePixelStream_s2mPipe_ready) begin
        readStage_counterOnePixelStream_rValid <= 1'b0;
      end
      if(readStage_counterOnePixelStream_s2mPipe_ready) begin
        readStage_counterOnePixelStream_s2mPipe_rValid <= readStage_counterOnePixelStream_s2mPipe_valid;
      end
      if(readStage_mainTwoPixelStream_valid) begin
        readStage_mainTwoPixelStream_rValid <= 1'b1;
      end
      if(readStage_mainTwoPixelStream_s2mPipe_ready) begin
        readStage_mainTwoPixelStream_rValid <= 1'b0;
      end
      if(readStage_mainTwoPixelStream_s2mPipe_ready) begin
        readStage_mainTwoPixelStream_s2mPipe_rValid <= readStage_mainTwoPixelStream_s2mPipe_valid;
      end
      if(readStage_counterTwoPixelStream_valid) begin
        readStage_counterTwoPixelStream_rValid <= 1'b1;
      end
      if(readStage_counterTwoPixelStream_s2mPipe_ready) begin
        readStage_counterTwoPixelStream_rValid <= 1'b0;
      end
      if(readStage_counterTwoPixelStream_s2mPipe_ready) begin
        readStage_counterTwoPixelStream_s2mPipe_rValid <= readStage_counterTwoPixelStream_s2mPipe_valid;
      end
      if(readStage_mainThreePixelStream_valid) begin
        readStage_mainThreePixelStream_rValid <= 1'b1;
      end
      if(readStage_mainThreePixelStream_s2mPipe_ready) begin
        readStage_mainThreePixelStream_rValid <= 1'b0;
      end
      if(readStage_mainThreePixelStream_s2mPipe_ready) begin
        readStage_mainThreePixelStream_s2mPipe_rValid <= readStage_mainThreePixelStream_s2mPipe_valid;
      end
      if(readStage_counterThreePixelStream_valid) begin
        readStage_counterThreePixelStream_rValid <= 1'b1;
      end
      if(readStage_counterThreePixelStream_s2mPipe_ready) begin
        readStage_counterThreePixelStream_rValid <= 1'b0;
      end
      if(readStage_counterThreePixelStream_s2mPipe_ready) begin
        readStage_counterThreePixelStream_s2mPipe_rValid <= readStage_counterThreePixelStream_s2mPipe_valid;
      end
      if(readStage_mainOneValidStream_valid) begin
        readStage_mainOneValidStream_rValid <= 1'b1;
      end
      if(readStage_mainOneValidStream_s2mPipe_ready) begin
        readStage_mainOneValidStream_rValid <= 1'b0;
      end
      if(readStage_mainOneValidStream_s2mPipe_ready) begin
        readStage_mainOneValidStream_s2mPipe_rValid <= readStage_mainOneValidStream_s2mPipe_valid;
      end
      if(readStage_counterOneValidStream_valid) begin
        readStage_counterOneValidStream_rValid <= 1'b1;
      end
      if(readStage_counterOneValidStream_s2mPipe_ready) begin
        readStage_counterOneValidStream_rValid <= 1'b0;
      end
      if(readStage_counterOneValidStream_s2mPipe_ready) begin
        readStage_counterOneValidStream_s2mPipe_rValid <= readStage_counterOneValidStream_s2mPipe_valid;
      end
      if(readStage_mainTwoValidStream_valid) begin
        readStage_mainTwoValidStream_rValid <= 1'b1;
      end
      if(readStage_mainTwoValidStream_s2mPipe_ready) begin
        readStage_mainTwoValidStream_rValid <= 1'b0;
      end
      if(readStage_mainTwoValidStream_s2mPipe_ready) begin
        readStage_mainTwoValidStream_s2mPipe_rValid <= readStage_mainTwoValidStream_s2mPipe_valid;
      end
      if(readStage_counterTwoValidStream_valid) begin
        readStage_counterTwoValidStream_rValid <= 1'b1;
      end
      if(readStage_counterTwoValidStream_s2mPipe_ready) begin
        readStage_counterTwoValidStream_rValid <= 1'b0;
      end
      if(readStage_counterTwoValidStream_s2mPipe_ready) begin
        readStage_counterTwoValidStream_s2mPipe_rValid <= readStage_counterTwoValidStream_s2mPipe_valid;
      end
      if(readStage_mainThreeValidStream_valid) begin
        readStage_mainThreeValidStream_rValid <= 1'b1;
      end
      if(readStage_mainThreeValidStream_s2mPipe_ready) begin
        readStage_mainThreeValidStream_rValid <= 1'b0;
      end
      if(readStage_mainThreeValidStream_s2mPipe_ready) begin
        readStage_mainThreeValidStream_s2mPipe_rValid <= readStage_mainThreeValidStream_s2mPipe_valid;
      end
      if(readStage_counterThreeValidStream_valid) begin
        readStage_counterThreeValidStream_rValid <= 1'b1;
      end
      if(readStage_counterThreeValidStream_s2mPipe_ready) begin
        readStage_counterThreeValidStream_rValid <= 1'b0;
      end
      if(readStage_counterThreeValidStream_s2mPipe_ready) begin
        readStage_counterThreeValidStream_s2mPipe_rValid <= readStage_counterThreeValidStream_s2mPipe_valid;
      end
      if(readStage_controlPipe_translated_valid) begin
        readStage_controlPipe_translated_rValid <= 1'b1;
      end
      if(readStage_controlPipe_translated_s2mPipe_ready) begin
        readStage_controlPipe_translated_rValid <= 1'b0;
      end
      if(readStage_controlPipe_translated_s2mPipe_ready) begin
        readStage_controlPipe_translated_s2mPipe_rValid <= readStage_controlPipe_translated_s2mPipe_valid;
      end
      if(compareStage_mainOnePixelStream_valid) begin
        compareStage_mainOnePixelStream_rValid <= 1'b1;
      end
      if(compareStage_mainOnePixelStream_s2mPipe_ready) begin
        compareStage_mainOnePixelStream_rValid <= 1'b0;
      end
      if(compareStage_mainOnePixelStream_s2mPipe_ready) begin
        compareStage_mainOnePixelStream_s2mPipe_rValid <= compareStage_mainOnePixelStream_s2mPipe_valid;
      end
      if(compareStage_counterOnePixelStream_valid) begin
        compareStage_counterOnePixelStream_rValid <= 1'b1;
      end
      if(compareStage_counterOnePixelStream_s2mPipe_ready) begin
        compareStage_counterOnePixelStream_rValid <= 1'b0;
      end
      if(compareStage_counterOnePixelStream_s2mPipe_ready) begin
        compareStage_counterOnePixelStream_s2mPipe_rValid <= compareStage_counterOnePixelStream_s2mPipe_valid;
      end
      if(compareStage_mainTwoPixelStream_valid) begin
        compareStage_mainTwoPixelStream_rValid <= 1'b1;
      end
      if(compareStage_mainTwoPixelStream_s2mPipe_ready) begin
        compareStage_mainTwoPixelStream_rValid <= 1'b0;
      end
      if(compareStage_mainTwoPixelStream_s2mPipe_ready) begin
        compareStage_mainTwoPixelStream_s2mPipe_rValid <= compareStage_mainTwoPixelStream_s2mPipe_valid;
      end
      if(compareStage_counterTwoPixelStream_valid) begin
        compareStage_counterTwoPixelStream_rValid <= 1'b1;
      end
      if(compareStage_counterTwoPixelStream_s2mPipe_ready) begin
        compareStage_counterTwoPixelStream_rValid <= 1'b0;
      end
      if(compareStage_counterTwoPixelStream_s2mPipe_ready) begin
        compareStage_counterTwoPixelStream_s2mPipe_rValid <= compareStage_counterTwoPixelStream_s2mPipe_valid;
      end
      if(compareStage_mainThreePixelStream_valid) begin
        compareStage_mainThreePixelStream_rValid <= 1'b1;
      end
      if(compareStage_mainThreePixelStream_s2mPipe_ready) begin
        compareStage_mainThreePixelStream_rValid <= 1'b0;
      end
      if(compareStage_mainThreePixelStream_s2mPipe_ready) begin
        compareStage_mainThreePixelStream_s2mPipe_rValid <= compareStage_mainThreePixelStream_s2mPipe_valid;
      end
      if(compareStage_counterThreePixelStream_valid) begin
        compareStage_counterThreePixelStream_rValid <= 1'b1;
      end
      if(compareStage_counterThreePixelStream_s2mPipe_ready) begin
        compareStage_counterThreePixelStream_rValid <= 1'b0;
      end
      if(compareStage_counterThreePixelStream_s2mPipe_ready) begin
        compareStage_counterThreePixelStream_s2mPipe_rValid <= compareStage_counterThreePixelStream_s2mPipe_valid;
      end
      if(compareStage_mainOneValidStream_valid) begin
        compareStage_mainOneValidStream_rValid <= 1'b1;
      end
      if(compareStage_mainOneValidStream_s2mPipe_ready) begin
        compareStage_mainOneValidStream_rValid <= 1'b0;
      end
      if(compareStage_mainOneValidStream_s2mPipe_ready) begin
        compareStage_mainOneValidStream_s2mPipe_rValid <= compareStage_mainOneValidStream_s2mPipe_valid;
      end
      if(compareStage_counterOneValidStream_valid) begin
        compareStage_counterOneValidStream_rValid <= 1'b1;
      end
      if(compareStage_counterOneValidStream_s2mPipe_ready) begin
        compareStage_counterOneValidStream_rValid <= 1'b0;
      end
      if(compareStage_counterOneValidStream_s2mPipe_ready) begin
        compareStage_counterOneValidStream_s2mPipe_rValid <= compareStage_counterOneValidStream_s2mPipe_valid;
      end
      if(compareStage_mainTwoValidStream_valid) begin
        compareStage_mainTwoValidStream_rValid <= 1'b1;
      end
      if(compareStage_mainTwoValidStream_s2mPipe_ready) begin
        compareStage_mainTwoValidStream_rValid <= 1'b0;
      end
      if(compareStage_mainTwoValidStream_s2mPipe_ready) begin
        compareStage_mainTwoValidStream_s2mPipe_rValid <= compareStage_mainTwoValidStream_s2mPipe_valid;
      end
      if(compareStage_counterTwoValidStream_valid) begin
        compareStage_counterTwoValidStream_rValid <= 1'b1;
      end
      if(compareStage_counterTwoValidStream_s2mPipe_ready) begin
        compareStage_counterTwoValidStream_rValid <= 1'b0;
      end
      if(compareStage_counterTwoValidStream_s2mPipe_ready) begin
        compareStage_counterTwoValidStream_s2mPipe_rValid <= compareStage_counterTwoValidStream_s2mPipe_valid;
      end
      if(compareStage_mainThreeValidStream_valid) begin
        compareStage_mainThreeValidStream_rValid <= 1'b1;
      end
      if(compareStage_mainThreeValidStream_s2mPipe_ready) begin
        compareStage_mainThreeValidStream_rValid <= 1'b0;
      end
      if(compareStage_mainThreeValidStream_s2mPipe_ready) begin
        compareStage_mainThreeValidStream_s2mPipe_rValid <= compareStage_mainThreeValidStream_s2mPipe_valid;
      end
      if(compareStage_counterThreeValidStream_valid) begin
        compareStage_counterThreeValidStream_rValid <= 1'b1;
      end
      if(compareStage_counterThreeValidStream_s2mPipe_ready) begin
        compareStage_counterThreeValidStream_rValid <= 1'b0;
      end
      if(compareStage_counterThreeValidStream_s2mPipe_ready) begin
        compareStage_counterThreeValidStream_s2mPipe_rValid <= compareStage_counterThreeValidStream_s2mPipe_valid;
      end
      if(compareStage_controlPipe_translated_valid) begin
        compareStage_controlPipe_translated_rValid <= 1'b1;
      end
      if(compareStage_controlPipe_translated_s2mPipe_ready) begin
        compareStage_controlPipe_translated_rValid <= 1'b0;
      end
      if(compareStage_controlPipe_translated_s2mPipe_ready) begin
        compareStage_controlPipe_translated_s2mPipe_rValid <= compareStage_controlPipe_translated_s2mPipe_valid;
      end
      if(diffStage_mainOnePixelStream_valid) begin
        diffStage_mainOnePixelStream_rValid <= 1'b1;
      end
      if(diffStage_mainOnePixelStream_s2mPipe_ready) begin
        diffStage_mainOnePixelStream_rValid <= 1'b0;
      end
      if(diffStage_mainOnePixelStream_s2mPipe_ready) begin
        diffStage_mainOnePixelStream_s2mPipe_rValid <= diffStage_mainOnePixelStream_s2mPipe_valid;
      end
      if(diffStage_counterOnePixelStream_valid) begin
        diffStage_counterOnePixelStream_rValid <= 1'b1;
      end
      if(diffStage_counterOnePixelStream_s2mPipe_ready) begin
        diffStage_counterOnePixelStream_rValid <= 1'b0;
      end
      if(diffStage_counterOnePixelStream_s2mPipe_ready) begin
        diffStage_counterOnePixelStream_s2mPipe_rValid <= diffStage_counterOnePixelStream_s2mPipe_valid;
      end
      if(diffStage_mainTwoPixelStream_valid) begin
        diffStage_mainTwoPixelStream_rValid <= 1'b1;
      end
      if(diffStage_mainTwoPixelStream_s2mPipe_ready) begin
        diffStage_mainTwoPixelStream_rValid <= 1'b0;
      end
      if(diffStage_mainTwoPixelStream_s2mPipe_ready) begin
        diffStage_mainTwoPixelStream_s2mPipe_rValid <= diffStage_mainTwoPixelStream_s2mPipe_valid;
      end
      if(diffStage_counterTwoPixelStream_valid) begin
        diffStage_counterTwoPixelStream_rValid <= 1'b1;
      end
      if(diffStage_counterTwoPixelStream_s2mPipe_ready) begin
        diffStage_counterTwoPixelStream_rValid <= 1'b0;
      end
      if(diffStage_counterTwoPixelStream_s2mPipe_ready) begin
        diffStage_counterTwoPixelStream_s2mPipe_rValid <= diffStage_counterTwoPixelStream_s2mPipe_valid;
      end
      if(diffStage_mainThreePixelStream_valid) begin
        diffStage_mainThreePixelStream_rValid <= 1'b1;
      end
      if(diffStage_mainThreePixelStream_s2mPipe_ready) begin
        diffStage_mainThreePixelStream_rValid <= 1'b0;
      end
      if(diffStage_mainThreePixelStream_s2mPipe_ready) begin
        diffStage_mainThreePixelStream_s2mPipe_rValid <= diffStage_mainThreePixelStream_s2mPipe_valid;
      end
      if(diffStage_counterThreePixelStream_valid) begin
        diffStage_counterThreePixelStream_rValid <= 1'b1;
      end
      if(diffStage_counterThreePixelStream_s2mPipe_ready) begin
        diffStage_counterThreePixelStream_rValid <= 1'b0;
      end
      if(diffStage_counterThreePixelStream_s2mPipe_ready) begin
        diffStage_counterThreePixelStream_s2mPipe_rValid <= diffStage_counterThreePixelStream_s2mPipe_valid;
      end
      if(diffStage_mainOneValidStream_valid) begin
        diffStage_mainOneValidStream_rValid <= 1'b1;
      end
      if(diffStage_mainOneValidStream_s2mPipe_ready) begin
        diffStage_mainOneValidStream_rValid <= 1'b0;
      end
      if(diffStage_mainOneValidStream_s2mPipe_ready) begin
        diffStage_mainOneValidStream_s2mPipe_rValid <= diffStage_mainOneValidStream_s2mPipe_valid;
      end
      if(diffStage_counterOneValidStream_valid) begin
        diffStage_counterOneValidStream_rValid <= 1'b1;
      end
      if(diffStage_counterOneValidStream_s2mPipe_ready) begin
        diffStage_counterOneValidStream_rValid <= 1'b0;
      end
      if(diffStage_counterOneValidStream_s2mPipe_ready) begin
        diffStage_counterOneValidStream_s2mPipe_rValid <= diffStage_counterOneValidStream_s2mPipe_valid;
      end
      if(diffStage_mainTwoValidStream_valid) begin
        diffStage_mainTwoValidStream_rValid <= 1'b1;
      end
      if(diffStage_mainTwoValidStream_s2mPipe_ready) begin
        diffStage_mainTwoValidStream_rValid <= 1'b0;
      end
      if(diffStage_mainTwoValidStream_s2mPipe_ready) begin
        diffStage_mainTwoValidStream_s2mPipe_rValid <= diffStage_mainTwoValidStream_s2mPipe_valid;
      end
      if(diffStage_counterTwoValidStream_valid) begin
        diffStage_counterTwoValidStream_rValid <= 1'b1;
      end
      if(diffStage_counterTwoValidStream_s2mPipe_ready) begin
        diffStage_counterTwoValidStream_rValid <= 1'b0;
      end
      if(diffStage_counterTwoValidStream_s2mPipe_ready) begin
        diffStage_counterTwoValidStream_s2mPipe_rValid <= diffStage_counterTwoValidStream_s2mPipe_valid;
      end
      if(diffStage_mainThreeValidStream_valid) begin
        diffStage_mainThreeValidStream_rValid <= 1'b1;
      end
      if(diffStage_mainThreeValidStream_s2mPipe_ready) begin
        diffStage_mainThreeValidStream_rValid <= 1'b0;
      end
      if(diffStage_mainThreeValidStream_s2mPipe_ready) begin
        diffStage_mainThreeValidStream_s2mPipe_rValid <= diffStage_mainThreeValidStream_s2mPipe_valid;
      end
      if(diffStage_counterThreeValidStream_valid) begin
        diffStage_counterThreeValidStream_rValid <= 1'b1;
      end
      if(diffStage_counterThreeValidStream_s2mPipe_ready) begin
        diffStage_counterThreeValidStream_rValid <= 1'b0;
      end
      if(diffStage_counterThreeValidStream_s2mPipe_ready) begin
        diffStage_counterThreeValidStream_s2mPipe_rValid <= diffStage_counterThreeValidStream_s2mPipe_valid;
      end
      if(resultStage_controlPipeBeforePipe_valid) begin
        resultStage_controlPipeBeforePipe_rValid <= 1'b1;
      end
      if(resultStage_controlPipeBeforePipe_s2mPipe_ready) begin
        resultStage_controlPipeBeforePipe_rValid <= 1'b0;
      end
      if(resultStage_controlPipeBeforePipe_s2mPipe_ready) begin
        resultStage_controlPipeBeforePipe_s2mPipe_rValid <= resultStage_controlPipeBeforePipe_s2mPipe_valid;
      end
      if(resultStage_pixelStream_valid) begin
        resultStage_pixelStream_rValid <= 1'b1;
      end
      if(resultStage_pixelStream_s2mPipe_ready) begin
        resultStage_pixelStream_rValid <= 1'b0;
      end
      if(resultStage_pixelStream_s2mPipe_ready) begin
        resultStage_pixelStream_s2mPipe_rValid <= resultStage_pixelStream_s2mPipe_valid;
      end
      if(when_SuperResolutionPart3_l1115) begin
        isHorizontalDirection <= resultStage_controlPipeBeforePipe_payload_isHorizontalMin;
        minDiff <= resultStage_controlPipeBeforePipe_payload_minDiff;
        candidatePixel <= resultStage_pixelStream_payload;
      end
      if(diffStage_controlPipe_fire) begin
        inValidMinDiff <= diffStage_controlPipe_payload_inValidMinDiff;
      end
      if(pixelsStream_valid) begin
        pixelsStream_rValid <= 1'b1;
      end
      if(pixelsStream_s2mPipe_ready) begin
        pixelsStream_rValid <= 1'b0;
      end
      if(pixelsStream_s2mPipe_ready) begin
        pixelsStream_s2mPipe_rValid <= pixelsStream_s2mPipe_valid;
      end
      controlStateMachine_stateReg <= controlStateMachine_stateNext;
      case(controlStateMachine_stateReg)
        controlStateMachine_enumDef_2_HOLD : begin
        end
        controlStateMachine_enumDef_2_PASS : begin
        end
        controlStateMachine_enumDef_2_EXTRA : begin
          if(when_SuperResolutionPart3_l1220) begin
            frameStart <= 1'b0;
          end
          if(when_SuperResolutionPart3_l1223) begin
            outReachRowEnd <= 1'b1;
          end
          if(when_SuperResolutionPart3_l1224) begin
            outReachFinalRow <= 1'b1;
          end
          if(when_SuperResolutionPart3_l1226) begin
            if(outReachFinalRow) begin
              startRead <= 1'b0;
              readDone <= 1'b1;
              outReachRowEnd <= 1'b0;
              outReachFinalRow <= 1'b0;
            end else begin
              outReachRowEnd <= 1'b0;
            end
          end
          if(controlStream_fire_6) begin
            if(outReachRowEnd) begin
              outReachRowEnd <= 1'b0;
            end
          end
          if(when_SuperResolutionPart3_l1247) begin
            if(when_SuperResolutionPart3_l1248) begin
              holdBuffer <= 1'b0;
            end
            if(when_SuperResolutionPart3_l1250) begin
              currentRowBuffer <= 2'b00;
            end else begin
              currentRowBuffer <= (currentRowBuffer + 2'b01);
            end
            if(when_SuperResolutionPart3_l1252) begin
              nextRowBuffer <= 2'b00;
            end else begin
              nextRowBuffer <= (nextRowBuffer + 2'b01);
            end
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(posedge clk) begin
    startIn_regNext <= startIn;
    startIn_regNext_1 <= startIn;
    if(pixelsIn_ready) begin
      pixelsIn_rData_pixel <= pixelsIn_payload_pixel;
      pixelsIn_rData_frameStart <= pixelsIn_payload_frameStart;
      pixelsIn_rData_rowEnd <= pixelsIn_payload_rowEnd;
      pixelsIn_rData_inpValid <= pixelsIn_payload_inpValid;
    end
    if(pixelsIn_s2mPipe_ready) begin
      pixelsIn_s2mPipe_rData_pixel <= pixelsIn_s2mPipe_payload_pixel;
      pixelsIn_s2mPipe_rData_frameStart <= pixelsIn_s2mPipe_payload_frameStart;
      pixelsIn_s2mPipe_rData_rowEnd <= pixelsIn_s2mPipe_payload_rowEnd;
      pixelsIn_s2mPipe_rData_inpValid <= pixelsIn_s2mPipe_payload_inpValid;
    end
    if(mainPixelAddrOneStream_ready) begin
      mainPixelAddrOneStream_rData <= mainPixelAddrOneStream_payload;
    end
    if(mainPixelAddrOneStream_s2mPipe_ready) begin
      mainPixelAddrOneStream_s2mPipe_rData <= mainPixelAddrOneStream_s2mPipe_payload;
    end
    if(CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_mainOnePixelStream_payload_1 <= CICC1851_readStage_mainOnePixelStream_payload;
    end
    if(CICC1851_1) begin
      CICC1851_readStage_mainOnePixelStream_payload_2 <= (CICC1851_mainPixelAddrOneStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_mainOnePixelStream_payload_1 : CICC1851_readStage_mainOnePixelStream_payload);
    end
    if(counterPixelAddrOneStream_ready) begin
      counterPixelAddrOneStream_rData <= counterPixelAddrOneStream_payload;
    end
    if(counterPixelAddrOneStream_s2mPipe_ready) begin
      counterPixelAddrOneStream_s2mPipe_rData <= counterPixelAddrOneStream_s2mPipe_payload;
    end
    if(CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_counterOnePixelStream_payload_1 <= CICC1851_readStage_counterOnePixelStream_payload;
    end
    if(CICC1851_2) begin
      CICC1851_readStage_counterOnePixelStream_payload_2 <= (CICC1851_counterPixelAddrOneStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_counterOnePixelStream_payload_1 : CICC1851_readStage_counterOnePixelStream_payload);
    end
    if(mainPixelAddrTwoStream_ready) begin
      mainPixelAddrTwoStream_rData <= mainPixelAddrTwoStream_payload;
    end
    if(mainPixelAddrTwoStream_s2mPipe_ready) begin
      mainPixelAddrTwoStream_s2mPipe_rData <= mainPixelAddrTwoStream_s2mPipe_payload;
    end
    if(CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_mainTwoPixelStream_payload_1 <= CICC1851_readStage_mainTwoPixelStream_payload;
    end
    if(CICC1851_3) begin
      CICC1851_readStage_mainTwoPixelStream_payload_2 <= (CICC1851_mainPixelAddrTwoStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_mainTwoPixelStream_payload_1 : CICC1851_readStage_mainTwoPixelStream_payload);
    end
    if(counterPixelAddrTwoStream_ready) begin
      counterPixelAddrTwoStream_rData <= counterPixelAddrTwoStream_payload;
    end
    if(counterPixelAddrTwoStream_s2mPipe_ready) begin
      counterPixelAddrTwoStream_s2mPipe_rData <= counterPixelAddrTwoStream_s2mPipe_payload;
    end
    if(CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_counterTwoPixelStream_payload_1 <= CICC1851_readStage_counterTwoPixelStream_payload;
    end
    if(CICC1851_4) begin
      CICC1851_readStage_counterTwoPixelStream_payload_2 <= (CICC1851_counterPixelAddrTwoStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_counterTwoPixelStream_payload_1 : CICC1851_readStage_counterTwoPixelStream_payload);
    end
    if(mainPixelAddrThreeStream_ready) begin
      mainPixelAddrThreeStream_rData <= mainPixelAddrThreeStream_payload;
    end
    if(mainPixelAddrThreeStream_s2mPipe_ready) begin
      mainPixelAddrThreeStream_s2mPipe_rData <= mainPixelAddrThreeStream_s2mPipe_payload;
    end
    if(CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_mainThreePixelStream_payload_1 <= CICC1851_readStage_mainThreePixelStream_payload;
    end
    if(CICC1851_5) begin
      CICC1851_readStage_mainThreePixelStream_payload_2 <= (CICC1851_mainPixelAddrThreeStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_mainThreePixelStream_payload_1 : CICC1851_readStage_mainThreePixelStream_payload);
    end
    if(counterPixelAddrThreeStream_ready) begin
      counterPixelAddrThreeStream_rData <= counterPixelAddrThreeStream_payload;
    end
    if(counterPixelAddrThreeStream_s2mPipe_ready) begin
      counterPixelAddrThreeStream_s2mPipe_rData <= counterPixelAddrThreeStream_s2mPipe_payload;
    end
    if(CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_counterThreePixelStream_payload_1 <= CICC1851_readStage_counterThreePixelStream_payload;
    end
    if(CICC1851_6) begin
      CICC1851_readStage_counterThreePixelStream_payload_2 <= (CICC1851_counterPixelAddrThreeStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_counterThreePixelStream_payload_1 : CICC1851_readStage_counterThreePixelStream_payload);
    end
    if(mainValidAddrOneStream_ready) begin
      mainValidAddrOneStream_rData <= mainValidAddrOneStream_payload;
    end
    if(mainValidAddrOneStream_s2mPipe_ready) begin
      mainValidAddrOneStream_s2mPipe_rData <= mainValidAddrOneStream_s2mPipe_payload;
    end
    if(CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_mainOneValidStream_payload_1 <= CICC1851_readStage_mainOneValidStream_payload;
    end
    if(CICC1851_7) begin
      CICC1851_readStage_mainOneValidStream_payload_2 <= (CICC1851_mainValidAddrOneStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_mainOneValidStream_payload_1 : CICC1851_readStage_mainOneValidStream_payload);
    end
    if(counterValidAddrOneStream_ready) begin
      counterValidAddrOneStream_rData <= counterValidAddrOneStream_payload;
    end
    if(counterValidAddrOneStream_s2mPipe_ready) begin
      counterValidAddrOneStream_s2mPipe_rData <= counterValidAddrOneStream_s2mPipe_payload;
    end
    if(CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_counterOneValidStream_payload_1 <= CICC1851_readStage_counterOneValidStream_payload;
    end
    if(CICC1851_8) begin
      CICC1851_readStage_counterOneValidStream_payload_2 <= (CICC1851_counterValidAddrOneStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_counterOneValidStream_payload_1 : CICC1851_readStage_counterOneValidStream_payload);
    end
    if(mainValidAddrTwoStream_ready) begin
      mainValidAddrTwoStream_rData <= mainValidAddrTwoStream_payload;
    end
    if(mainValidAddrTwoStream_s2mPipe_ready) begin
      mainValidAddrTwoStream_s2mPipe_rData <= mainValidAddrTwoStream_s2mPipe_payload;
    end
    if(CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_mainTwoValidStream_payload_1 <= CICC1851_readStage_mainTwoValidStream_payload;
    end
    if(CICC1851_9) begin
      CICC1851_readStage_mainTwoValidStream_payload_2 <= (CICC1851_mainValidAddrTwoStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_mainTwoValidStream_payload_1 : CICC1851_readStage_mainTwoValidStream_payload);
    end
    if(counterValidAddrTwoStream_ready) begin
      counterValidAddrTwoStream_rData <= counterValidAddrTwoStream_payload;
    end
    if(counterValidAddrTwoStream_s2mPipe_ready) begin
      counterValidAddrTwoStream_s2mPipe_rData <= counterValidAddrTwoStream_s2mPipe_payload;
    end
    if(CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_counterTwoValidStream_payload_1 <= CICC1851_readStage_counterTwoValidStream_payload;
    end
    if(CICC1851_10) begin
      CICC1851_readStage_counterTwoValidStream_payload_2 <= (CICC1851_counterValidAddrTwoStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_counterTwoValidStream_payload_1 : CICC1851_readStage_counterTwoValidStream_payload);
    end
    if(mainValidAddrThreeStream_ready) begin
      mainValidAddrThreeStream_rData <= mainValidAddrThreeStream_payload;
    end
    if(mainValidAddrThreeStream_s2mPipe_ready) begin
      mainValidAddrThreeStream_s2mPipe_rData <= mainValidAddrThreeStream_s2mPipe_payload;
    end
    if(CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_mainThreeValidStream_payload_1 <= CICC1851_readStage_mainThreeValidStream_payload;
    end
    if(CICC1851_11) begin
      CICC1851_readStage_mainThreeValidStream_payload_2 <= (CICC1851_mainValidAddrThreeStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_mainThreeValidStream_payload_1 : CICC1851_readStage_mainThreeValidStream_payload);
    end
    if(counterValidAddrThreeStream_ready) begin
      counterValidAddrThreeStream_rData <= counterValidAddrThreeStream_payload;
    end
    if(counterValidAddrThreeStream_s2mPipe_ready) begin
      counterValidAddrThreeStream_s2mPipe_rData <= counterValidAddrThreeStream_s2mPipe_payload;
    end
    if(CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_counterThreeValidStream_payload_1 <= CICC1851_readStage_counterThreeValidStream_payload;
    end
    if(CICC1851_12) begin
      CICC1851_readStage_counterThreeValidStream_payload_2 <= (CICC1851_counterValidAddrThreeStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_counterThreeValidStream_payload_1 : CICC1851_readStage_counterThreeValidStream_payload);
    end
    if(controlStream_ready) begin
      controlStream_rData_frameStart <= controlStream_payload_frameStart;
      controlStream_rData_rowEnd <= controlStream_payload_rowEnd;
      controlStream_rData_pipeValid <= controlStream_payload_pipeValid;
      controlStream_rData_firstRow <= controlStream_payload_firstRow;
      controlStream_rData_lastRow <= controlStream_payload_lastRow;
      controlStream_rData_finalResult <= controlStream_payload_finalResult;
      controlStream_rData_mainCompare <= controlStream_payload_mainCompare;
      controlStream_rData_counterCompare <= controlStream_payload_counterCompare;
      controlStream_rData_horizontalCompare <= controlStream_payload_horizontalCompare;
      controlStream_rData_verticalCompare <= controlStream_payload_verticalCompare;
      controlStream_rData_mainDiff <= controlStream_payload_mainDiff;
      controlStream_rData_counterDiff <= controlStream_payload_counterDiff;
      controlStream_rData_horizontalDiff <= controlStream_payload_horizontalDiff;
      controlStream_rData_verticalDiff <= controlStream_payload_verticalDiff;
      controlStream_rData_isHorizontalMin <= controlStream_payload_isHorizontalMin;
      controlStream_rData_minDiff <= controlStream_payload_minDiff;
      controlStream_rData_currentPosition <= controlStream_payload_currentPosition;
      controlStream_rData_nextPosition <= controlStream_payload_nextPosition;
      controlStream_rData_horizontalDirectionValid <= controlStream_payload_horizontalDirectionValid;
      controlStream_rData_verticalDirectionValid <= controlStream_payload_verticalDirectionValid;
      controlStream_rData_mainDirectionValid <= controlStream_payload_mainDirectionValid;
      controlStream_rData_counterDirectionValid <= controlStream_payload_counterDirectionValid;
      controlStream_rData_inValidMinDiff <= controlStream_payload_inValidMinDiff;
    end
    if(controlStream_s2mPipe_ready) begin
      controlStream_s2mPipe_rData_frameStart <= controlStream_s2mPipe_payload_frameStart;
      controlStream_s2mPipe_rData_rowEnd <= controlStream_s2mPipe_payload_rowEnd;
      controlStream_s2mPipe_rData_pipeValid <= controlStream_s2mPipe_payload_pipeValid;
      controlStream_s2mPipe_rData_firstRow <= controlStream_s2mPipe_payload_firstRow;
      controlStream_s2mPipe_rData_lastRow <= controlStream_s2mPipe_payload_lastRow;
      controlStream_s2mPipe_rData_finalResult <= controlStream_s2mPipe_payload_finalResult;
      controlStream_s2mPipe_rData_mainCompare <= controlStream_s2mPipe_payload_mainCompare;
      controlStream_s2mPipe_rData_counterCompare <= controlStream_s2mPipe_payload_counterCompare;
      controlStream_s2mPipe_rData_horizontalCompare <= controlStream_s2mPipe_payload_horizontalCompare;
      controlStream_s2mPipe_rData_verticalCompare <= controlStream_s2mPipe_payload_verticalCompare;
      controlStream_s2mPipe_rData_mainDiff <= controlStream_s2mPipe_payload_mainDiff;
      controlStream_s2mPipe_rData_counterDiff <= controlStream_s2mPipe_payload_counterDiff;
      controlStream_s2mPipe_rData_horizontalDiff <= controlStream_s2mPipe_payload_horizontalDiff;
      controlStream_s2mPipe_rData_verticalDiff <= controlStream_s2mPipe_payload_verticalDiff;
      controlStream_s2mPipe_rData_isHorizontalMin <= controlStream_s2mPipe_payload_isHorizontalMin;
      controlStream_s2mPipe_rData_minDiff <= controlStream_s2mPipe_payload_minDiff;
      controlStream_s2mPipe_rData_currentPosition <= controlStream_s2mPipe_payload_currentPosition;
      controlStream_s2mPipe_rData_nextPosition <= controlStream_s2mPipe_payload_nextPosition;
      controlStream_s2mPipe_rData_horizontalDirectionValid <= controlStream_s2mPipe_payload_horizontalDirectionValid;
      controlStream_s2mPipe_rData_verticalDirectionValid <= controlStream_s2mPipe_payload_verticalDirectionValid;
      controlStream_s2mPipe_rData_mainDirectionValid <= controlStream_s2mPipe_payload_mainDirectionValid;
      controlStream_s2mPipe_rData_counterDirectionValid <= controlStream_s2mPipe_payload_counterDirectionValid;
      controlStream_s2mPipe_rData_inValidMinDiff <= controlStream_s2mPipe_payload_inValidMinDiff;
    end
    if(controlStream_s2mPipe_m2sPipe_ready) begin
      controlStream_s2mPipe_m2sPipe_rData_frameStart <= controlStream_s2mPipe_m2sPipe_payload_frameStart;
      controlStream_s2mPipe_m2sPipe_rData_rowEnd <= controlStream_s2mPipe_m2sPipe_payload_rowEnd;
      controlStream_s2mPipe_m2sPipe_rData_pipeValid <= controlStream_s2mPipe_m2sPipe_payload_pipeValid;
      controlStream_s2mPipe_m2sPipe_rData_firstRow <= controlStream_s2mPipe_m2sPipe_payload_firstRow;
      controlStream_s2mPipe_m2sPipe_rData_lastRow <= controlStream_s2mPipe_m2sPipe_payload_lastRow;
      controlStream_s2mPipe_m2sPipe_rData_finalResult <= controlStream_s2mPipe_m2sPipe_payload_finalResult;
      controlStream_s2mPipe_m2sPipe_rData_mainCompare <= controlStream_s2mPipe_m2sPipe_payload_mainCompare;
      controlStream_s2mPipe_m2sPipe_rData_counterCompare <= controlStream_s2mPipe_m2sPipe_payload_counterCompare;
      controlStream_s2mPipe_m2sPipe_rData_horizontalCompare <= controlStream_s2mPipe_m2sPipe_payload_horizontalCompare;
      controlStream_s2mPipe_m2sPipe_rData_verticalCompare <= controlStream_s2mPipe_m2sPipe_payload_verticalCompare;
      controlStream_s2mPipe_m2sPipe_rData_mainDiff <= controlStream_s2mPipe_m2sPipe_payload_mainDiff;
      controlStream_s2mPipe_m2sPipe_rData_counterDiff <= controlStream_s2mPipe_m2sPipe_payload_counterDiff;
      controlStream_s2mPipe_m2sPipe_rData_horizontalDiff <= controlStream_s2mPipe_m2sPipe_payload_horizontalDiff;
      controlStream_s2mPipe_m2sPipe_rData_verticalDiff <= controlStream_s2mPipe_m2sPipe_payload_verticalDiff;
      controlStream_s2mPipe_m2sPipe_rData_isHorizontalMin <= controlStream_s2mPipe_m2sPipe_payload_isHorizontalMin;
      controlStream_s2mPipe_m2sPipe_rData_minDiff <= controlStream_s2mPipe_m2sPipe_payload_minDiff;
      controlStream_s2mPipe_m2sPipe_rData_currentPosition <= controlStream_s2mPipe_m2sPipe_payload_currentPosition;
      controlStream_s2mPipe_m2sPipe_rData_nextPosition <= controlStream_s2mPipe_m2sPipe_payload_nextPosition;
      controlStream_s2mPipe_m2sPipe_rData_horizontalDirectionValid <= controlStream_s2mPipe_m2sPipe_payload_horizontalDirectionValid;
      controlStream_s2mPipe_m2sPipe_rData_verticalDirectionValid <= controlStream_s2mPipe_m2sPipe_payload_verticalDirectionValid;
      controlStream_s2mPipe_m2sPipe_rData_mainDirectionValid <= controlStream_s2mPipe_m2sPipe_payload_mainDirectionValid;
      controlStream_s2mPipe_m2sPipe_rData_counterDirectionValid <= controlStream_s2mPipe_m2sPipe_payload_counterDirectionValid;
      controlStream_s2mPipe_m2sPipe_rData_inValidMinDiff <= controlStream_s2mPipe_m2sPipe_payload_inValidMinDiff;
    end
    if(controlStream_s2mPipe_m2sPipe_m2sPipe_ready) begin
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_frameStart <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_frameStart;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_rowEnd <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_rowEnd;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_pipeValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_pipeValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_firstRow <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_firstRow;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_lastRow <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_lastRow;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_finalResult <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_finalResult;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_horizontalCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_horizontalCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_verticalCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_verticalCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_horizontalDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_horizontalDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_verticalDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_verticalDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_isHorizontalMin <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_isHorizontalMin;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_minDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_minDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_currentPosition <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_currentPosition;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_nextPosition <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_nextPosition;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_horizontalDirectionValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_horizontalDirectionValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_verticalDirectionValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_verticalDirectionValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainDirectionValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDirectionValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterDirectionValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDirectionValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_inValidMinDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_inValidMinDiff;
    end
    if(controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready) begin
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_frameStart <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_frameStart;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_rowEnd <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_rowEnd;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_pipeValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_pipeValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_firstRow <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_firstRow;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_lastRow <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_lastRow;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_finalResult <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_finalResult;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_horizontalCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_horizontalCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_verticalCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_verticalCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_horizontalDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_horizontalDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_verticalDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_verticalDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_isHorizontalMin <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_isHorizontalMin;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_minDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_minDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_currentPosition <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_currentPosition;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_nextPosition <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_nextPosition;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_horizontalDirectionValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_horizontalDirectionValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_verticalDirectionValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_verticalDirectionValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainDirectionValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainDirectionValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterDirectionValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterDirectionValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_inValidMinDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_inValidMinDiff;
    end
    if(readStage_mainOnePixelStream_ready) begin
      readStage_mainOnePixelStream_rData <= readStage_mainOnePixelStream_payload;
    end
    if(readStage_mainOnePixelStream_s2mPipe_ready) begin
      readStage_mainOnePixelStream_s2mPipe_rData <= readStage_mainOnePixelStream_s2mPipe_payload;
    end
    if(readStage_counterOnePixelStream_ready) begin
      readStage_counterOnePixelStream_rData <= readStage_counterOnePixelStream_payload;
    end
    if(readStage_counterOnePixelStream_s2mPipe_ready) begin
      readStage_counterOnePixelStream_s2mPipe_rData <= readStage_counterOnePixelStream_s2mPipe_payload;
    end
    if(readStage_mainTwoPixelStream_ready) begin
      readStage_mainTwoPixelStream_rData <= readStage_mainTwoPixelStream_payload;
    end
    if(readStage_mainTwoPixelStream_s2mPipe_ready) begin
      readStage_mainTwoPixelStream_s2mPipe_rData <= readStage_mainTwoPixelStream_s2mPipe_payload;
    end
    if(readStage_counterTwoPixelStream_ready) begin
      readStage_counterTwoPixelStream_rData <= readStage_counterTwoPixelStream_payload;
    end
    if(readStage_counterTwoPixelStream_s2mPipe_ready) begin
      readStage_counterTwoPixelStream_s2mPipe_rData <= readStage_counterTwoPixelStream_s2mPipe_payload;
    end
    if(readStage_mainThreePixelStream_ready) begin
      readStage_mainThreePixelStream_rData <= readStage_mainThreePixelStream_payload;
    end
    if(readStage_mainThreePixelStream_s2mPipe_ready) begin
      readStage_mainThreePixelStream_s2mPipe_rData <= readStage_mainThreePixelStream_s2mPipe_payload;
    end
    if(readStage_counterThreePixelStream_ready) begin
      readStage_counterThreePixelStream_rData <= readStage_counterThreePixelStream_payload;
    end
    if(readStage_counterThreePixelStream_s2mPipe_ready) begin
      readStage_counterThreePixelStream_s2mPipe_rData <= readStage_counterThreePixelStream_s2mPipe_payload;
    end
    if(readStage_mainOneValidStream_ready) begin
      readStage_mainOneValidStream_rData <= readStage_mainOneValidStream_payload;
    end
    if(readStage_mainOneValidStream_s2mPipe_ready) begin
      readStage_mainOneValidStream_s2mPipe_rData <= readStage_mainOneValidStream_s2mPipe_payload;
    end
    if(readStage_counterOneValidStream_ready) begin
      readStage_counterOneValidStream_rData <= readStage_counterOneValidStream_payload;
    end
    if(readStage_counterOneValidStream_s2mPipe_ready) begin
      readStage_counterOneValidStream_s2mPipe_rData <= readStage_counterOneValidStream_s2mPipe_payload;
    end
    if(readStage_mainTwoValidStream_ready) begin
      readStage_mainTwoValidStream_rData <= readStage_mainTwoValidStream_payload;
    end
    if(readStage_mainTwoValidStream_s2mPipe_ready) begin
      readStage_mainTwoValidStream_s2mPipe_rData <= readStage_mainTwoValidStream_s2mPipe_payload;
    end
    if(readStage_counterTwoValidStream_ready) begin
      readStage_counterTwoValidStream_rData <= readStage_counterTwoValidStream_payload;
    end
    if(readStage_counterTwoValidStream_s2mPipe_ready) begin
      readStage_counterTwoValidStream_s2mPipe_rData <= readStage_counterTwoValidStream_s2mPipe_payload;
    end
    if(readStage_mainThreeValidStream_ready) begin
      readStage_mainThreeValidStream_rData <= readStage_mainThreeValidStream_payload;
    end
    if(readStage_mainThreeValidStream_s2mPipe_ready) begin
      readStage_mainThreeValidStream_s2mPipe_rData <= readStage_mainThreeValidStream_s2mPipe_payload;
    end
    if(readStage_counterThreeValidStream_ready) begin
      readStage_counterThreeValidStream_rData <= readStage_counterThreeValidStream_payload;
    end
    if(readStage_counterThreeValidStream_s2mPipe_ready) begin
      readStage_counterThreeValidStream_s2mPipe_rData <= readStage_counterThreeValidStream_s2mPipe_payload;
    end
    if(readStage_controlPipe_translated_ready) begin
      readStage_controlPipe_translated_rData_frameStart <= readStage_controlPipe_translated_payload_frameStart;
      readStage_controlPipe_translated_rData_rowEnd <= readStage_controlPipe_translated_payload_rowEnd;
      readStage_controlPipe_translated_rData_pipeValid <= readStage_controlPipe_translated_payload_pipeValid;
      readStage_controlPipe_translated_rData_firstRow <= readStage_controlPipe_translated_payload_firstRow;
      readStage_controlPipe_translated_rData_lastRow <= readStage_controlPipe_translated_payload_lastRow;
      readStage_controlPipe_translated_rData_finalResult <= readStage_controlPipe_translated_payload_finalResult;
      readStage_controlPipe_translated_rData_mainCompare <= readStage_controlPipe_translated_payload_mainCompare;
      readStage_controlPipe_translated_rData_counterCompare <= readStage_controlPipe_translated_payload_counterCompare;
      readStage_controlPipe_translated_rData_horizontalCompare <= readStage_controlPipe_translated_payload_horizontalCompare;
      readStage_controlPipe_translated_rData_verticalCompare <= readStage_controlPipe_translated_payload_verticalCompare;
      readStage_controlPipe_translated_rData_mainDiff <= readStage_controlPipe_translated_payload_mainDiff;
      readStage_controlPipe_translated_rData_counterDiff <= readStage_controlPipe_translated_payload_counterDiff;
      readStage_controlPipe_translated_rData_horizontalDiff <= readStage_controlPipe_translated_payload_horizontalDiff;
      readStage_controlPipe_translated_rData_verticalDiff <= readStage_controlPipe_translated_payload_verticalDiff;
      readStage_controlPipe_translated_rData_isHorizontalMin <= readStage_controlPipe_translated_payload_isHorizontalMin;
      readStage_controlPipe_translated_rData_minDiff <= readStage_controlPipe_translated_payload_minDiff;
      readStage_controlPipe_translated_rData_currentPosition <= readStage_controlPipe_translated_payload_currentPosition;
      readStage_controlPipe_translated_rData_nextPosition <= readStage_controlPipe_translated_payload_nextPosition;
      readStage_controlPipe_translated_rData_horizontalDirectionValid <= readStage_controlPipe_translated_payload_horizontalDirectionValid;
      readStage_controlPipe_translated_rData_verticalDirectionValid <= readStage_controlPipe_translated_payload_verticalDirectionValid;
      readStage_controlPipe_translated_rData_mainDirectionValid <= readStage_controlPipe_translated_payload_mainDirectionValid;
      readStage_controlPipe_translated_rData_counterDirectionValid <= readStage_controlPipe_translated_payload_counterDirectionValid;
      readStage_controlPipe_translated_rData_inValidMinDiff <= readStage_controlPipe_translated_payload_inValidMinDiff;
    end
    if(readStage_controlPipe_translated_s2mPipe_ready) begin
      readStage_controlPipe_translated_s2mPipe_rData_frameStart <= readStage_controlPipe_translated_s2mPipe_payload_frameStart;
      readStage_controlPipe_translated_s2mPipe_rData_rowEnd <= readStage_controlPipe_translated_s2mPipe_payload_rowEnd;
      readStage_controlPipe_translated_s2mPipe_rData_pipeValid <= readStage_controlPipe_translated_s2mPipe_payload_pipeValid;
      readStage_controlPipe_translated_s2mPipe_rData_firstRow <= readStage_controlPipe_translated_s2mPipe_payload_firstRow;
      readStage_controlPipe_translated_s2mPipe_rData_lastRow <= readStage_controlPipe_translated_s2mPipe_payload_lastRow;
      readStage_controlPipe_translated_s2mPipe_rData_finalResult <= readStage_controlPipe_translated_s2mPipe_payload_finalResult;
      readStage_controlPipe_translated_s2mPipe_rData_mainCompare <= readStage_controlPipe_translated_s2mPipe_payload_mainCompare;
      readStage_controlPipe_translated_s2mPipe_rData_counterCompare <= readStage_controlPipe_translated_s2mPipe_payload_counterCompare;
      readStage_controlPipe_translated_s2mPipe_rData_horizontalCompare <= readStage_controlPipe_translated_s2mPipe_payload_horizontalCompare;
      readStage_controlPipe_translated_s2mPipe_rData_verticalCompare <= readStage_controlPipe_translated_s2mPipe_payload_verticalCompare;
      readStage_controlPipe_translated_s2mPipe_rData_mainDiff <= readStage_controlPipe_translated_s2mPipe_payload_mainDiff;
      readStage_controlPipe_translated_s2mPipe_rData_counterDiff <= readStage_controlPipe_translated_s2mPipe_payload_counterDiff;
      readStage_controlPipe_translated_s2mPipe_rData_horizontalDiff <= readStage_controlPipe_translated_s2mPipe_payload_horizontalDiff;
      readStage_controlPipe_translated_s2mPipe_rData_verticalDiff <= readStage_controlPipe_translated_s2mPipe_payload_verticalDiff;
      readStage_controlPipe_translated_s2mPipe_rData_isHorizontalMin <= readStage_controlPipe_translated_s2mPipe_payload_isHorizontalMin;
      readStage_controlPipe_translated_s2mPipe_rData_minDiff <= readStage_controlPipe_translated_s2mPipe_payload_minDiff;
      readStage_controlPipe_translated_s2mPipe_rData_currentPosition <= readStage_controlPipe_translated_s2mPipe_payload_currentPosition;
      readStage_controlPipe_translated_s2mPipe_rData_nextPosition <= readStage_controlPipe_translated_s2mPipe_payload_nextPosition;
      readStage_controlPipe_translated_s2mPipe_rData_horizontalDirectionValid <= readStage_controlPipe_translated_s2mPipe_payload_horizontalDirectionValid;
      readStage_controlPipe_translated_s2mPipe_rData_verticalDirectionValid <= readStage_controlPipe_translated_s2mPipe_payload_verticalDirectionValid;
      readStage_controlPipe_translated_s2mPipe_rData_mainDirectionValid <= readStage_controlPipe_translated_s2mPipe_payload_mainDirectionValid;
      readStage_controlPipe_translated_s2mPipe_rData_counterDirectionValid <= readStage_controlPipe_translated_s2mPipe_payload_counterDirectionValid;
      readStage_controlPipe_translated_s2mPipe_rData_inValidMinDiff <= readStage_controlPipe_translated_s2mPipe_payload_inValidMinDiff;
    end
    if(compareStage_mainOnePixelStream_ready) begin
      compareStage_mainOnePixelStream_rData <= compareStage_mainOnePixelStream_payload;
    end
    if(compareStage_mainOnePixelStream_s2mPipe_ready) begin
      compareStage_mainOnePixelStream_s2mPipe_rData <= compareStage_mainOnePixelStream_s2mPipe_payload;
    end
    if(compareStage_counterOnePixelStream_ready) begin
      compareStage_counterOnePixelStream_rData <= compareStage_counterOnePixelStream_payload;
    end
    if(compareStage_counterOnePixelStream_s2mPipe_ready) begin
      compareStage_counterOnePixelStream_s2mPipe_rData <= compareStage_counterOnePixelStream_s2mPipe_payload;
    end
    if(compareStage_mainTwoPixelStream_ready) begin
      compareStage_mainTwoPixelStream_rData <= compareStage_mainTwoPixelStream_payload;
    end
    if(compareStage_mainTwoPixelStream_s2mPipe_ready) begin
      compareStage_mainTwoPixelStream_s2mPipe_rData <= compareStage_mainTwoPixelStream_s2mPipe_payload;
    end
    if(compareStage_counterTwoPixelStream_ready) begin
      compareStage_counterTwoPixelStream_rData <= compareStage_counterTwoPixelStream_payload;
    end
    if(compareStage_counterTwoPixelStream_s2mPipe_ready) begin
      compareStage_counterTwoPixelStream_s2mPipe_rData <= compareStage_counterTwoPixelStream_s2mPipe_payload;
    end
    if(compareStage_mainThreePixelStream_ready) begin
      compareStage_mainThreePixelStream_rData <= compareStage_mainThreePixelStream_payload;
    end
    if(compareStage_mainThreePixelStream_s2mPipe_ready) begin
      compareStage_mainThreePixelStream_s2mPipe_rData <= compareStage_mainThreePixelStream_s2mPipe_payload;
    end
    if(compareStage_counterThreePixelStream_ready) begin
      compareStage_counterThreePixelStream_rData <= compareStage_counterThreePixelStream_payload;
    end
    if(compareStage_counterThreePixelStream_s2mPipe_ready) begin
      compareStage_counterThreePixelStream_s2mPipe_rData <= compareStage_counterThreePixelStream_s2mPipe_payload;
    end
    if(compareStage_mainOneValidStream_ready) begin
      compareStage_mainOneValidStream_rData <= compareStage_mainOneValidStream_payload;
    end
    if(compareStage_mainOneValidStream_s2mPipe_ready) begin
      compareStage_mainOneValidStream_s2mPipe_rData <= compareStage_mainOneValidStream_s2mPipe_payload;
    end
    if(compareStage_counterOneValidStream_ready) begin
      compareStage_counterOneValidStream_rData <= compareStage_counterOneValidStream_payload;
    end
    if(compareStage_counterOneValidStream_s2mPipe_ready) begin
      compareStage_counterOneValidStream_s2mPipe_rData <= compareStage_counterOneValidStream_s2mPipe_payload;
    end
    if(compareStage_mainTwoValidStream_ready) begin
      compareStage_mainTwoValidStream_rData <= compareStage_mainTwoValidStream_payload;
    end
    if(compareStage_mainTwoValidStream_s2mPipe_ready) begin
      compareStage_mainTwoValidStream_s2mPipe_rData <= compareStage_mainTwoValidStream_s2mPipe_payload;
    end
    if(compareStage_counterTwoValidStream_ready) begin
      compareStage_counterTwoValidStream_rData <= compareStage_counterTwoValidStream_payload;
    end
    if(compareStage_counterTwoValidStream_s2mPipe_ready) begin
      compareStage_counterTwoValidStream_s2mPipe_rData <= compareStage_counterTwoValidStream_s2mPipe_payload;
    end
    if(compareStage_mainThreeValidStream_ready) begin
      compareStage_mainThreeValidStream_rData <= compareStage_mainThreeValidStream_payload;
    end
    if(compareStage_mainThreeValidStream_s2mPipe_ready) begin
      compareStage_mainThreeValidStream_s2mPipe_rData <= compareStage_mainThreeValidStream_s2mPipe_payload;
    end
    if(compareStage_counterThreeValidStream_ready) begin
      compareStage_counterThreeValidStream_rData <= compareStage_counterThreeValidStream_payload;
    end
    if(compareStage_counterThreeValidStream_s2mPipe_ready) begin
      compareStage_counterThreeValidStream_s2mPipe_rData <= compareStage_counterThreeValidStream_s2mPipe_payload;
    end
    if(compareStage_controlPipe_translated_ready) begin
      compareStage_controlPipe_translated_rData_frameStart <= compareStage_controlPipe_translated_payload_frameStart;
      compareStage_controlPipe_translated_rData_rowEnd <= compareStage_controlPipe_translated_payload_rowEnd;
      compareStage_controlPipe_translated_rData_pipeValid <= compareStage_controlPipe_translated_payload_pipeValid;
      compareStage_controlPipe_translated_rData_firstRow <= compareStage_controlPipe_translated_payload_firstRow;
      compareStage_controlPipe_translated_rData_lastRow <= compareStage_controlPipe_translated_payload_lastRow;
      compareStage_controlPipe_translated_rData_finalResult <= compareStage_controlPipe_translated_payload_finalResult;
      compareStage_controlPipe_translated_rData_mainCompare <= compareStage_controlPipe_translated_payload_mainCompare;
      compareStage_controlPipe_translated_rData_counterCompare <= compareStage_controlPipe_translated_payload_counterCompare;
      compareStage_controlPipe_translated_rData_horizontalCompare <= compareStage_controlPipe_translated_payload_horizontalCompare;
      compareStage_controlPipe_translated_rData_verticalCompare <= compareStage_controlPipe_translated_payload_verticalCompare;
      compareStage_controlPipe_translated_rData_mainDiff <= compareStage_controlPipe_translated_payload_mainDiff;
      compareStage_controlPipe_translated_rData_counterDiff <= compareStage_controlPipe_translated_payload_counterDiff;
      compareStage_controlPipe_translated_rData_horizontalDiff <= compareStage_controlPipe_translated_payload_horizontalDiff;
      compareStage_controlPipe_translated_rData_verticalDiff <= compareStage_controlPipe_translated_payload_verticalDiff;
      compareStage_controlPipe_translated_rData_isHorizontalMin <= compareStage_controlPipe_translated_payload_isHorizontalMin;
      compareStage_controlPipe_translated_rData_minDiff <= compareStage_controlPipe_translated_payload_minDiff;
      compareStage_controlPipe_translated_rData_currentPosition <= compareStage_controlPipe_translated_payload_currentPosition;
      compareStage_controlPipe_translated_rData_nextPosition <= compareStage_controlPipe_translated_payload_nextPosition;
      compareStage_controlPipe_translated_rData_horizontalDirectionValid <= compareStage_controlPipe_translated_payload_horizontalDirectionValid;
      compareStage_controlPipe_translated_rData_verticalDirectionValid <= compareStage_controlPipe_translated_payload_verticalDirectionValid;
      compareStage_controlPipe_translated_rData_mainDirectionValid <= compareStage_controlPipe_translated_payload_mainDirectionValid;
      compareStage_controlPipe_translated_rData_counterDirectionValid <= compareStage_controlPipe_translated_payload_counterDirectionValid;
      compareStage_controlPipe_translated_rData_inValidMinDiff <= compareStage_controlPipe_translated_payload_inValidMinDiff;
    end
    if(compareStage_controlPipe_translated_s2mPipe_ready) begin
      compareStage_controlPipe_translated_s2mPipe_rData_frameStart <= compareStage_controlPipe_translated_s2mPipe_payload_frameStart;
      compareStage_controlPipe_translated_s2mPipe_rData_rowEnd <= compareStage_controlPipe_translated_s2mPipe_payload_rowEnd;
      compareStage_controlPipe_translated_s2mPipe_rData_pipeValid <= compareStage_controlPipe_translated_s2mPipe_payload_pipeValid;
      compareStage_controlPipe_translated_s2mPipe_rData_firstRow <= compareStage_controlPipe_translated_s2mPipe_payload_firstRow;
      compareStage_controlPipe_translated_s2mPipe_rData_lastRow <= compareStage_controlPipe_translated_s2mPipe_payload_lastRow;
      compareStage_controlPipe_translated_s2mPipe_rData_finalResult <= compareStage_controlPipe_translated_s2mPipe_payload_finalResult;
      compareStage_controlPipe_translated_s2mPipe_rData_mainCompare <= compareStage_controlPipe_translated_s2mPipe_payload_mainCompare;
      compareStage_controlPipe_translated_s2mPipe_rData_counterCompare <= compareStage_controlPipe_translated_s2mPipe_payload_counterCompare;
      compareStage_controlPipe_translated_s2mPipe_rData_horizontalCompare <= compareStage_controlPipe_translated_s2mPipe_payload_horizontalCompare;
      compareStage_controlPipe_translated_s2mPipe_rData_verticalCompare <= compareStage_controlPipe_translated_s2mPipe_payload_verticalCompare;
      compareStage_controlPipe_translated_s2mPipe_rData_mainDiff <= compareStage_controlPipe_translated_s2mPipe_payload_mainDiff;
      compareStage_controlPipe_translated_s2mPipe_rData_counterDiff <= compareStage_controlPipe_translated_s2mPipe_payload_counterDiff;
      compareStage_controlPipe_translated_s2mPipe_rData_horizontalDiff <= compareStage_controlPipe_translated_s2mPipe_payload_horizontalDiff;
      compareStage_controlPipe_translated_s2mPipe_rData_verticalDiff <= compareStage_controlPipe_translated_s2mPipe_payload_verticalDiff;
      compareStage_controlPipe_translated_s2mPipe_rData_isHorizontalMin <= compareStage_controlPipe_translated_s2mPipe_payload_isHorizontalMin;
      compareStage_controlPipe_translated_s2mPipe_rData_minDiff <= compareStage_controlPipe_translated_s2mPipe_payload_minDiff;
      compareStage_controlPipe_translated_s2mPipe_rData_currentPosition <= compareStage_controlPipe_translated_s2mPipe_payload_currentPosition;
      compareStage_controlPipe_translated_s2mPipe_rData_nextPosition <= compareStage_controlPipe_translated_s2mPipe_payload_nextPosition;
      compareStage_controlPipe_translated_s2mPipe_rData_horizontalDirectionValid <= compareStage_controlPipe_translated_s2mPipe_payload_horizontalDirectionValid;
      compareStage_controlPipe_translated_s2mPipe_rData_verticalDirectionValid <= compareStage_controlPipe_translated_s2mPipe_payload_verticalDirectionValid;
      compareStage_controlPipe_translated_s2mPipe_rData_mainDirectionValid <= compareStage_controlPipe_translated_s2mPipe_payload_mainDirectionValid;
      compareStage_controlPipe_translated_s2mPipe_rData_counterDirectionValid <= compareStage_controlPipe_translated_s2mPipe_payload_counterDirectionValid;
      compareStage_controlPipe_translated_s2mPipe_rData_inValidMinDiff <= compareStage_controlPipe_translated_s2mPipe_payload_inValidMinDiff;
    end
    if(diffStage_mainOnePixelStream_ready) begin
      diffStage_mainOnePixelStream_rData <= diffStage_mainOnePixelStream_payload;
    end
    if(diffStage_mainOnePixelStream_s2mPipe_ready) begin
      diffStage_mainOnePixelStream_s2mPipe_rData <= diffStage_mainOnePixelStream_s2mPipe_payload;
    end
    if(diffStage_counterOnePixelStream_ready) begin
      diffStage_counterOnePixelStream_rData <= diffStage_counterOnePixelStream_payload;
    end
    if(diffStage_counterOnePixelStream_s2mPipe_ready) begin
      diffStage_counterOnePixelStream_s2mPipe_rData <= diffStage_counterOnePixelStream_s2mPipe_payload;
    end
    if(diffStage_mainTwoPixelStream_ready) begin
      diffStage_mainTwoPixelStream_rData <= diffStage_mainTwoPixelStream_payload;
    end
    if(diffStage_mainTwoPixelStream_s2mPipe_ready) begin
      diffStage_mainTwoPixelStream_s2mPipe_rData <= diffStage_mainTwoPixelStream_s2mPipe_payload;
    end
    if(diffStage_counterTwoPixelStream_ready) begin
      diffStage_counterTwoPixelStream_rData <= diffStage_counterTwoPixelStream_payload;
    end
    if(diffStage_counterTwoPixelStream_s2mPipe_ready) begin
      diffStage_counterTwoPixelStream_s2mPipe_rData <= diffStage_counterTwoPixelStream_s2mPipe_payload;
    end
    if(diffStage_mainThreePixelStream_ready) begin
      diffStage_mainThreePixelStream_rData <= diffStage_mainThreePixelStream_payload;
    end
    if(diffStage_mainThreePixelStream_s2mPipe_ready) begin
      diffStage_mainThreePixelStream_s2mPipe_rData <= diffStage_mainThreePixelStream_s2mPipe_payload;
    end
    if(diffStage_counterThreePixelStream_ready) begin
      diffStage_counterThreePixelStream_rData <= diffStage_counterThreePixelStream_payload;
    end
    if(diffStage_counterThreePixelStream_s2mPipe_ready) begin
      diffStage_counterThreePixelStream_s2mPipe_rData <= diffStage_counterThreePixelStream_s2mPipe_payload;
    end
    if(diffStage_mainOneValidStream_ready) begin
      diffStage_mainOneValidStream_rData <= diffStage_mainOneValidStream_payload;
    end
    if(diffStage_mainOneValidStream_s2mPipe_ready) begin
      diffStage_mainOneValidStream_s2mPipe_rData <= diffStage_mainOneValidStream_s2mPipe_payload;
    end
    if(diffStage_counterOneValidStream_ready) begin
      diffStage_counterOneValidStream_rData <= diffStage_counterOneValidStream_payload;
    end
    if(diffStage_counterOneValidStream_s2mPipe_ready) begin
      diffStage_counterOneValidStream_s2mPipe_rData <= diffStage_counterOneValidStream_s2mPipe_payload;
    end
    if(diffStage_mainTwoValidStream_ready) begin
      diffStage_mainTwoValidStream_rData <= diffStage_mainTwoValidStream_payload;
    end
    if(diffStage_mainTwoValidStream_s2mPipe_ready) begin
      diffStage_mainTwoValidStream_s2mPipe_rData <= diffStage_mainTwoValidStream_s2mPipe_payload;
    end
    if(diffStage_counterTwoValidStream_ready) begin
      diffStage_counterTwoValidStream_rData <= diffStage_counterTwoValidStream_payload;
    end
    if(diffStage_counterTwoValidStream_s2mPipe_ready) begin
      diffStage_counterTwoValidStream_s2mPipe_rData <= diffStage_counterTwoValidStream_s2mPipe_payload;
    end
    if(diffStage_mainThreeValidStream_ready) begin
      diffStage_mainThreeValidStream_rData <= diffStage_mainThreeValidStream_payload;
    end
    if(diffStage_mainThreeValidStream_s2mPipe_ready) begin
      diffStage_mainThreeValidStream_s2mPipe_rData <= diffStage_mainThreeValidStream_s2mPipe_payload;
    end
    if(diffStage_counterThreeValidStream_ready) begin
      diffStage_counterThreeValidStream_rData <= diffStage_counterThreeValidStream_payload;
    end
    if(diffStage_counterThreeValidStream_s2mPipe_ready) begin
      diffStage_counterThreeValidStream_s2mPipe_rData <= diffStage_counterThreeValidStream_s2mPipe_payload;
    end
    if(resultStage_controlPipeBeforePipe_ready) begin
      resultStage_controlPipeBeforePipe_rData_frameStart <= resultStage_controlPipeBeforePipe_payload_frameStart;
      resultStage_controlPipeBeforePipe_rData_rowEnd <= resultStage_controlPipeBeforePipe_payload_rowEnd;
      resultStage_controlPipeBeforePipe_rData_pipeValid <= resultStage_controlPipeBeforePipe_payload_pipeValid;
      resultStage_controlPipeBeforePipe_rData_firstRow <= resultStage_controlPipeBeforePipe_payload_firstRow;
      resultStage_controlPipeBeforePipe_rData_lastRow <= resultStage_controlPipeBeforePipe_payload_lastRow;
      resultStage_controlPipeBeforePipe_rData_finalResult <= resultStage_controlPipeBeforePipe_payload_finalResult;
      resultStage_controlPipeBeforePipe_rData_mainCompare <= resultStage_controlPipeBeforePipe_payload_mainCompare;
      resultStage_controlPipeBeforePipe_rData_counterCompare <= resultStage_controlPipeBeforePipe_payload_counterCompare;
      resultStage_controlPipeBeforePipe_rData_horizontalCompare <= resultStage_controlPipeBeforePipe_payload_horizontalCompare;
      resultStage_controlPipeBeforePipe_rData_verticalCompare <= resultStage_controlPipeBeforePipe_payload_verticalCompare;
      resultStage_controlPipeBeforePipe_rData_mainDiff <= resultStage_controlPipeBeforePipe_payload_mainDiff;
      resultStage_controlPipeBeforePipe_rData_counterDiff <= resultStage_controlPipeBeforePipe_payload_counterDiff;
      resultStage_controlPipeBeforePipe_rData_horizontalDiff <= resultStage_controlPipeBeforePipe_payload_horizontalDiff;
      resultStage_controlPipeBeforePipe_rData_verticalDiff <= resultStage_controlPipeBeforePipe_payload_verticalDiff;
      resultStage_controlPipeBeforePipe_rData_isHorizontalMin <= resultStage_controlPipeBeforePipe_payload_isHorizontalMin;
      resultStage_controlPipeBeforePipe_rData_minDiff <= resultStage_controlPipeBeforePipe_payload_minDiff;
      resultStage_controlPipeBeforePipe_rData_currentPosition <= resultStage_controlPipeBeforePipe_payload_currentPosition;
      resultStage_controlPipeBeforePipe_rData_nextPosition <= resultStage_controlPipeBeforePipe_payload_nextPosition;
      resultStage_controlPipeBeforePipe_rData_horizontalDirectionValid <= resultStage_controlPipeBeforePipe_payload_horizontalDirectionValid;
      resultStage_controlPipeBeforePipe_rData_verticalDirectionValid <= resultStage_controlPipeBeforePipe_payload_verticalDirectionValid;
      resultStage_controlPipeBeforePipe_rData_mainDirectionValid <= resultStage_controlPipeBeforePipe_payload_mainDirectionValid;
      resultStage_controlPipeBeforePipe_rData_counterDirectionValid <= resultStage_controlPipeBeforePipe_payload_counterDirectionValid;
      resultStage_controlPipeBeforePipe_rData_inValidMinDiff <= resultStage_controlPipeBeforePipe_payload_inValidMinDiff;
    end
    if(resultStage_controlPipeBeforePipe_s2mPipe_ready) begin
      resultStage_controlPipeBeforePipe_s2mPipe_rData_frameStart <= resultStage_controlPipeBeforePipe_s2mPipe_payload_frameStart;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_rowEnd <= resultStage_controlPipeBeforePipe_s2mPipe_payload_rowEnd;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_pipeValid <= resultStage_controlPipeBeforePipe_s2mPipe_payload_pipeValid;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_firstRow <= resultStage_controlPipeBeforePipe_s2mPipe_payload_firstRow;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_lastRow <= resultStage_controlPipeBeforePipe_s2mPipe_payload_lastRow;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_finalResult <= resultStage_controlPipeBeforePipe_s2mPipe_payload_finalResult;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_mainCompare <= resultStage_controlPipeBeforePipe_s2mPipe_payload_mainCompare;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_counterCompare <= resultStage_controlPipeBeforePipe_s2mPipe_payload_counterCompare;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_horizontalCompare <= resultStage_controlPipeBeforePipe_s2mPipe_payload_horizontalCompare;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_verticalCompare <= resultStage_controlPipeBeforePipe_s2mPipe_payload_verticalCompare;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_mainDiff <= resultStage_controlPipeBeforePipe_s2mPipe_payload_mainDiff;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_counterDiff <= resultStage_controlPipeBeforePipe_s2mPipe_payload_counterDiff;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_horizontalDiff <= resultStage_controlPipeBeforePipe_s2mPipe_payload_horizontalDiff;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_verticalDiff <= resultStage_controlPipeBeforePipe_s2mPipe_payload_verticalDiff;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_isHorizontalMin <= resultStage_controlPipeBeforePipe_s2mPipe_payload_isHorizontalMin;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_minDiff <= resultStage_controlPipeBeforePipe_s2mPipe_payload_minDiff;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_currentPosition <= resultStage_controlPipeBeforePipe_s2mPipe_payload_currentPosition;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_nextPosition <= resultStage_controlPipeBeforePipe_s2mPipe_payload_nextPosition;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_horizontalDirectionValid <= resultStage_controlPipeBeforePipe_s2mPipe_payload_horizontalDirectionValid;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_verticalDirectionValid <= resultStage_controlPipeBeforePipe_s2mPipe_payload_verticalDirectionValid;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_mainDirectionValid <= resultStage_controlPipeBeforePipe_s2mPipe_payload_mainDirectionValid;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_counterDirectionValid <= resultStage_controlPipeBeforePipe_s2mPipe_payload_counterDirectionValid;
      resultStage_controlPipeBeforePipe_s2mPipe_rData_inValidMinDiff <= resultStage_controlPipeBeforePipe_s2mPipe_payload_inValidMinDiff;
    end
    if(resultStage_pixelStream_ready) begin
      resultStage_pixelStream_rData <= resultStage_pixelStream_payload;
    end
    if(resultStage_pixelStream_s2mPipe_ready) begin
      resultStage_pixelStream_s2mPipe_rData <= resultStage_pixelStream_s2mPipe_payload;
    end
    if(pixelsStream_ready) begin
      pixelsStream_rData_pixel <= pixelsStream_payload_pixel;
      pixelsStream_rData_frameStart <= pixelsStream_payload_frameStart;
      pixelsStream_rData_rowEnd <= pixelsStream_payload_rowEnd;
    end
    if(pixelsStream_s2mPipe_ready) begin
      pixelsStream_s2mPipe_rData_pixel <= pixelsStream_s2mPipe_payload_pixel;
      pixelsStream_s2mPipe_rData_frameStart <= pixelsStream_s2mPipe_payload_frameStart;
      pixelsStream_s2mPipe_rData_rowEnd <= pixelsStream_s2mPipe_payload_rowEnd;
    end
  end


endmodule

module SuperResolutionPart2 (
  input               pixelsIn_valid,
  output reg          pixelsIn_ready,
  input      [7:0]    pixelsIn_payload_pixel,
  input               pixelsIn_payload_frameStart,
  input               pixelsIn_payload_rowEnd,
  input               startIn,
  input               inpThreeDoneIn,
  output reg          pixelsOut_valid,
  input               pixelsOut_ready,
  output reg [7:0]    pixelsOut_payload_pixel,
  output reg          pixelsOut_payload_frameStart,
  output reg          pixelsOut_payload_rowEnd,
  output reg          pixelsOut_payload_inpValid,
  output reg          startOut,
  output reg          inpTwoDoneOut,
  input      [7:0]    thresholdIn,
  input      [9:0]    widthIn,
  input      [9:0]    heightIn,
  input               clk,
  input               resetn
);
  localparam controlStateMachine_enumDef_1_BOOT = 3'd0;
  localparam controlStateMachine_enumDef_1_HOLD = 3'd1;
  localparam controlStateMachine_enumDef_1_PASS = 3'd2;
  localparam controlStateMachine_enumDef_1_ONCE = 3'd3;
  localparam controlStateMachine_enumDef_1_TWICE = 3'd4;

  reg        [7:0]    CICC1851_lineBufferOne_port1;
  reg        [7:0]    CICC1851_lineBufferOne_port2;
  reg        [7:0]    CICC1851_lineBufferTwo_port1;
  reg        [7:0]    CICC1851_lineBufferTwo_port2;
  reg        [7:0]    CICC1851_lineBufferOdd_port1;
  wire                diffStage_controlPipe_fork_io_input_ready;
  wire                diffStage_controlPipe_fork_io_outputs_0_valid;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_frameStart;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_rowEnd;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_passMode;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_passValid;
  wire       [2:0]    diffStage_controlPipe_fork_io_outputs_0_payload_onceMode;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_onceValid;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_mainCompare;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_counterCompare;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_payload_mainDiff;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_payload_counterDiff;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_twiceCompValid;
  wire       [2:0]    diffStage_controlPipe_fork_io_outputs_0_payload_twiceMode;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_inpValidFlag;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_oddValid;
  wire                diffStage_controlPipe_fork_io_outputs_1_valid;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_frameStart;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_rowEnd;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_passMode;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_passValid;
  wire       [2:0]    diffStage_controlPipe_fork_io_outputs_1_payload_onceMode;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_onceValid;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_mainCompare;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_counterCompare;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_twiceCompValid;
  wire       [2:0]    diffStage_controlPipe_fork_io_outputs_1_payload_twiceMode;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_inpValidFlag;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_oddValid;
  wire       [10:0]   CICC1851_bufferRowCount_valueNext;
  wire       [0:0]    CICC1851_bufferRowCount_valueNext_1;
  wire       [10:0]   CICC1851_bufferWAddr_valueNext;
  wire       [0:0]    CICC1851_bufferWAddr_valueNext_1;
  wire       [11:0]   CICC1851_outPixelAddr_valueNext;
  wire       [0:0]    CICC1851_outPixelAddr_valueNext_1;
  wire       [11:0]   CICC1851_outRowCount_valueNext;
  wire       [0:0]    CICC1851_outRowCount_valueNext_1;
  wire       [11:0]   CICC1851_alreadySendRow_valueNext;
  wire       [0:0]    CICC1851_alreadySendRow_valueNext_1;
  wire       [11:0]   CICC1851_alreadySendCountInRow_valueNext;
  wire       [0:0]    CICC1851_alreadySendCountInRow_valueNext_1;
  wire       [11:0]   CICC1851_mainAddrOne;
  wire       [11:0]   CICC1851_counterAddrOne;
  wire       [11:0]   CICC1851_mainAddrTwo;
  wire       [11:0]   CICC1851_counterAddrTwo;
  wire       [11:0]   CICC1851_oddAddr;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l181;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l181_1;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l181_2;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l182;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l182_1;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l182_2;
  wire       [10:0]   CICC1851_when_SuperResolutionPart2_l195;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l218;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l234;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l234_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l234_2;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l235;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l235_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l235_2;
  wire       [7:0]    CICC1851_lineBufferOne_port;
  wire                CICC1851_lineBufferOne_port_1;
  wire       [7:0]    CICC1851_lineBufferOdd_port;
  wire                CICC1851_lineBufferOdd_port_1;
  wire       [7:0]    CICC1851_lineBufferTwo_port;
  wire                CICC1851_lineBufferTwo_port_1;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_1;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_2;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_3;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_4;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_5;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_6;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_7;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_8;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_9;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_10;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_11;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_12;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_13;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_14;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_15;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_16;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_17;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_18;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_19;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l763;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l763_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l763_2;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l764;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l764_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l764_2;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l783;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l785;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l787;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l789;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l793;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l796;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l799;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l802;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l560;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l560_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l602;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l602_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l602_2;
  wire       [2:0]    CICC1851_when_SuperResolutionPart2_l602_3;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l603;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l603_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l605;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l605_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l605_2;
  wire       [2:0]    CICC1851_when_SuperResolutionPart2_l605_3;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l606;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l606_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l606_2;
  wire       [1:0]    CICC1851_when_SuperResolutionPart2_l606_3;
  wire       [11:0]   CICC1851_when_SuperResolutionPart2_l609;
  wire       [11:0]   CICC1851_mainAddrOne_1;
  wire       [11:0]   CICC1851_mainAddrOne_2;
  wire       [11:0]   CICC1851_mainAddrTwo_1;
  wire       [11:0]   CICC1851_mainAddrTwo_2;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l667;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l667_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l667_2;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l667_3;
  wire       [1:0]    CICC1851_when_SuperResolutionPart2_l667_4;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l668;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l668_1;
  wire       [12:0]   CICC1851_when_SuperResolutionPart2_l668_2;
  wire       [1:0]    CICC1851_when_SuperResolutionPart2_l668_3;
  wire       [11:0]   CICC1851_mainAddrOne_3;
  wire       [11:0]   CICC1851_mainAddrOne_4;
  wire       [11:0]   CICC1851_mainAddrTwo_3;
  wire       [11:0]   CICC1851_mainAddrTwo_4;
  wire       [1:0]    CICC1851_controls_onceMode;
  wire       [1:0]    CICC1851_controls_onceMode_1;
  wire       [11:0]   CICC1851_mainAddrOne_5;
  wire       [11:0]   CICC1851_mainAddrOne_6;
  wire       [11:0]   CICC1851_counterAddrOne_1;
  wire       [11:0]   CICC1851_counterAddrOne_2;
  wire       [11:0]   CICC1851_counterAddrOne_3;
  wire       [11:0]   CICC1851_counterAddrOne_4;
  wire       [0:0]    CICC1851_controls_onceMode_2;
  wire       [11:0]   CICC1851_mainAddrTwo_5;
  wire       [11:0]   CICC1851_mainAddrTwo_6;
  wire       [11:0]   CICC1851_counterAddrTwo_1;
  wire       [11:0]   CICC1851_counterAddrTwo_2;
  wire       [11:0]   CICC1851_counterAddrTwo_3;
  wire       [11:0]   CICC1851_counterAddrTwo_4;
  wire       [11:0]   CICC1851_mainAddrOne_7;
  wire       [11:0]   CICC1851_mainAddrOne_8;
  wire       [11:0]   CICC1851_mainAddrOne_9;
  wire       [11:0]   CICC1851_mainAddrOne_10;
  wire       [12:0]   CICC1851_counterAddrOne_5;
  wire       [12:0]   CICC1851_counterAddrOne_6;
  wire       [12:0]   CICC1851_counterAddrOne_7;
  wire       [1:0]    CICC1851_counterAddrOne_8;
  wire       [1:0]    CICC1851_controls_twiceMode;
  wire       [11:0]   CICC1851_mainAddrTwo_7;
  wire       [11:0]   CICC1851_mainAddrTwo_8;
  wire       [1:0]    CICC1851_controls_twiceMode_1;
  wire       [11:0]   CICC1851_mainAddrTwo_9;
  wire       [11:0]   CICC1851_mainAddrTwo_10;
  wire       [12:0]   CICC1851_counterAddrTwo_5;
  wire       [12:0]   CICC1851_counterAddrTwo_6;
  wire       [12:0]   CICC1851_counterAddrTwo_7;
  wire       [1:0]    CICC1851_counterAddrTwo_8;
  wire       [11:0]   CICC1851_mainAddrOne_11;
  wire       [11:0]   CICC1851_mainAddrOne_12;
  wire       [11:0]   CICC1851_counterAddrTwo_9;
  wire       [11:0]   CICC1851_counterAddrTwo_10;
  wire       [11:0]   CICC1851_mainAddrTwo_11;
  wire       [11:0]   CICC1851_mainAddrTwo_12;
  wire       [11:0]   CICC1851_counterAddrOne_9;
  wire       [11:0]   CICC1851_counterAddrOne_10;
  wire       [12:0]   CICC1851_mainAddrTwo_13;
  wire       [12:0]   CICC1851_mainAddrTwo_14;
  wire       [12:0]   CICC1851_mainAddrTwo_15;
  wire       [1:0]    CICC1851_mainAddrTwo_16;
  wire       [12:0]   CICC1851_counterAddrOne_11;
  wire       [12:0]   CICC1851_counterAddrOne_12;
  wire       [12:0]   CICC1851_counterAddrOne_13;
  wire       [1:0]    CICC1851_counterAddrOne_14;
  wire       [0:0]    CICC1851_controls_twiceMode_2;
  wire       [11:0]   CICC1851_mainAddrTwo_17;
  wire       [11:0]   CICC1851_mainAddrTwo_18;
  wire       [11:0]   CICC1851_counterAddrOne_15;
  wire       [11:0]   CICC1851_counterAddrOne_16;
  wire       [11:0]   CICC1851_mainAddrOne_13;
  wire       [11:0]   CICC1851_mainAddrOne_14;
  wire       [11:0]   CICC1851_counterAddrTwo_11;
  wire       [11:0]   CICC1851_counterAddrTwo_12;
  wire       [12:0]   CICC1851_mainAddrOne_15;
  wire       [12:0]   CICC1851_mainAddrOne_16;
  wire       [12:0]   CICC1851_mainAddrOne_17;
  wire       [1:0]    CICC1851_mainAddrOne_18;
  wire       [12:0]   CICC1851_counterAddrTwo_13;
  wire       [12:0]   CICC1851_counterAddrTwo_14;
  wire       [12:0]   CICC1851_counterAddrTwo_15;
  wire       [1:0]    CICC1851_counterAddrTwo_16;
  reg                 inpTwoDone;
  reg                 startIn_regNext;
  wire                when_SuperResolutionPart2_l40;
  reg                 readDone;
  wire                when_SuperResolutionPart2_l43;
  reg                 startRead;
  wire                when_SuperResolutionPart2_l46;
  wire                when_SuperResolutionPart2_l46_1;
  reg                 slaveStart;
  wire                pixelsIn_fire;
  wire                when_SuperResolutionPart2_l49;
  wire                when_SuperResolutionPart2_l49_1;
  reg                 frameStart;
  reg        [7:0]    inpThreshold;
  reg        [9:0]    bmpWidth;
  reg        [9:0]    bmpHeight;
  reg                 holdBuffer;
  wire                when_SuperResolutionPart2_l64;
  reg                 writeDone;
  wire                when_SuperResolutionPart2_l67;
  reg                 bufferRowCount_willIncrement;
  reg                 bufferRowCount_willClear;
  reg        [10:0]   bufferRowCount_valueNext;
  reg        [10:0]   bufferRowCount_value;
  wire                bufferRowCount_willOverflowIfInc;
  wire                bufferRowCount_willOverflow;
  reg                 bufferReuse;
  reg                 bufferEnable;
  wire                when_SuperResolutionPart2_l76;
  wire                when_SuperResolutionPart2_l76_1;
  reg        [1:0]    bufferSwitch;
  reg                 nextRowBuffer;
  wire                when_SuperResolutionPart2_l82;
  reg                 bufferWAddr_willIncrement;
  reg                 bufferWAddr_willClear;
  reg        [10:0]   bufferWAddr_valueNext;
  reg        [10:0]   bufferWAddr_value;
  wire                bufferWAddr_willOverflowIfInc;
  wire                bufferWAddr_willOverflow;
  reg                 outPixelAddr_willIncrement;
  reg                 outPixelAddr_willClear;
  reg        [11:0]   outPixelAddr_valueNext;
  reg        [11:0]   outPixelAddr_value;
  wire                outPixelAddr_willOverflowIfInc;
  wire                outPixelAddr_willOverflow;
  reg                 outRowCount_willIncrement;
  reg                 outRowCount_willClear;
  reg        [11:0]   outRowCount_valueNext;
  reg        [11:0]   outRowCount_value;
  wire                outRowCount_willOverflowIfInc;
  wire                outRowCount_willOverflow;
  reg                 alreadySendRow_willIncrement;
  reg                 alreadySendRow_willClear;
  reg        [11:0]   alreadySendRow_valueNext;
  reg        [11:0]   alreadySendRow_value;
  wire                alreadySendRow_willOverflowIfInc;
  wire                alreadySendRow_willOverflow;
  reg                 alreadySendCountInRow_willIncrement;
  reg                 alreadySendCountInRow_willClear;
  reg        [11:0]   alreadySendCountInRow_valueNext;
  reg        [11:0]   alreadySendCountInRow_value;
  wire                alreadySendCountInRow_willOverflowIfInc;
  wire                alreadySendCountInRow_willOverflow;
  reg                 alreadyReachRowEnd;
  reg                 alreadyReachFinalRow;
  reg                 outReachRowEnd;
  reg                 outReachFinalRow;
  reg                 bufferReachRowEnd;
  reg                 bufferReachFinalRow;
  reg                 oddBufferRow;
  reg                 startIn_regNext_1;
  wire                when_SuperResolutionPart2_l106;
  reg                 zeroInFourOutPixelAddr;
  reg                 startIn_regNext_2;
  wire                when_SuperResolutionPart2_l108;
  reg                 oneInFourOutPixelAddr;
  reg                 startIn_regNext_3;
  wire                when_SuperResolutionPart2_l109;
  reg                 twoInFourOutPixelAddr;
  reg                 startIn_regNext_4;
  wire                when_SuperResolutionPart2_l110;
  reg                 threeInFourOutPixelAddr;
  reg                 startIn_regNext_5;
  wire                when_SuperResolutionPart2_l111;
  reg                 zeroInFourOutRow;
  reg                 startIn_regNext_6;
  wire                when_SuperResolutionPart2_l113;
  reg                 oneInFourOutRow;
  reg                 startIn_regNext_7;
  wire                when_SuperResolutionPart2_l114;
  reg                 twoInFourOutRow;
  reg                 startIn_regNext_8;
  wire                when_SuperResolutionPart2_l115;
  reg                 threeInFourOutRow;
  reg                 startIn_regNext_9;
  wire                when_SuperResolutionPart2_l116;
  wire       [2:0]    currentState;
  reg                 willHoldToTwice;
  reg                 startIn_regNext_10;
  wire                when_SuperResolutionPart2_l120;
  reg                 willPassToHoldCaseOne;
  reg                 startIn_regNext_11;
  wire                when_SuperResolutionPart2_l121;
  reg                 willPassToHoldCaseTwo;
  reg                 startIn_regNext_12;
  wire                when_SuperResolutionPart2_l122;
  reg                 holdWillPassToHoldCaseTwo;
  reg                 startIn_regNext_13;
  wire                when_SuperResolutionPart2_l123;
  reg                 willOnceToHoldCaseOne;
  reg                 startIn_regNext_14;
  wire                when_SuperResolutionPart2_l124;
  reg                 willOnceToHoldCaseTwo;
  reg                 startIn_regNext_15;
  wire                when_SuperResolutionPart2_l125;
  reg                 willOnceToHoldCaseThree;
  reg                 startIn_regNext_16;
  wire                when_SuperResolutionPart2_l126;
  wire                when_SuperResolutionPart2_l134;
  reg        [10:0]   mainAddrOne;
  reg        [10:0]   counterAddrOne;
  reg        [10:0]   mainAddrTwo;
  reg        [10:0]   counterAddrTwo;
  wire       [10:0]   oddAddr;
  wire                validStream_valid;
  reg                 validStream_ready;
  wire                controlStream_valid;
  wire                controlStream_ready;
  wire                controlStream_payload_frameStart;
  wire                controlStream_payload_rowEnd;
  wire                controlStream_payload_passMode;
  wire                controlStream_payload_passValid;
  wire       [2:0]    controlStream_payload_onceMode;
  wire                controlStream_payload_onceValid;
  wire                controlStream_payload_mainCompare;
  wire                controlStream_payload_counterCompare;
  wire       [7:0]    controlStream_payload_mainDiff;
  wire       [7:0]    controlStream_payload_counterDiff;
  wire                controlStream_payload_twiceCompValid;
  wire       [2:0]    controlStream_payload_twiceMode;
  wire                controlStream_payload_inpValidFlag;
  wire                controlStream_payload_oddValid;
  reg                 controls_frameStart;
  reg                 controls_rowEnd;
  reg                 controls_passMode;
  reg                 controls_passValid;
  reg        [2:0]    controls_onceMode;
  reg                 controls_onceValid;
  wire                controls_mainCompare;
  wire                controls_counterCompare;
  wire       [7:0]    controls_mainDiff;
  wire       [7:0]    controls_counterDiff;
  reg                 controls_twiceCompValid;
  reg        [2:0]    controls_twiceMode;
  reg                 controls_inpValidFlag;
  reg                 controls_oddValid;
  wire       [31:0]   CICC1851_controls_frameStart;
  wire                mainAddrOneStream_valid;
  wire                mainAddrOneStream_ready;
  wire       [10:0]   mainAddrOneStream_payload;
  wire                counterAddrOneStream_valid;
  wire                counterAddrOneStream_ready;
  wire       [10:0]   counterAddrOneStream_payload;
  wire                mainAddrTwoStream_valid;
  wire                mainAddrTwoStream_ready;
  wire       [10:0]   mainAddrTwoStream_payload;
  wire                counterAddrTwoStream_valid;
  wire                counterAddrTwoStream_ready;
  wire       [10:0]   counterAddrTwoStream_payload;
  wire                oddAddrStream_valid;
  wire                oddAddrStream_ready;
  wire       [10:0]   oddAddrStream_payload;
  wire                pixelsIn_s2mPipe_valid;
  reg                 pixelsIn_s2mPipe_ready;
  wire       [7:0]    pixelsIn_s2mPipe_payload_pixel;
  wire                pixelsIn_s2mPipe_payload_frameStart;
  wire                pixelsIn_s2mPipe_payload_rowEnd;
  reg                 pixelsIn_rValid;
  reg        [7:0]    pixelsIn_rData_pixel;
  reg                 pixelsIn_rData_frameStart;
  reg                 pixelsIn_rData_rowEnd;
  wire                pixelsIn_s2mPipe_m2sPipe_valid;
  wire                pixelsIn_s2mPipe_m2sPipe_ready;
  wire       [7:0]    pixelsIn_s2mPipe_m2sPipe_payload_pixel;
  wire                pixelsIn_s2mPipe_m2sPipe_payload_frameStart;
  wire                pixelsIn_s2mPipe_m2sPipe_payload_rowEnd;
  reg                 pixelsIn_s2mPipe_rValid;
  reg        [7:0]    pixelsIn_s2mPipe_rData_pixel;
  reg                 pixelsIn_s2mPipe_rData_frameStart;
  reg                 pixelsIn_s2mPipe_rData_rowEnd;
  wire                when_Stream_l368;
  wire                passPixels_valid;
  wire                passPixels_ready;
  wire       [7:0]    passPixels_payload_pixel;
  wire                passPixels_payload_frameStart;
  wire                passPixels_payload_rowEnd;
  wire                passPixels_fire;
  wire                when_SuperResolutionPart2_l181;
  wire                passPixels_fire_1;
  wire                when_SuperResolutionPart2_l182;
  wire                passPixels_fire_2;
  wire                when_SuperResolutionPart2_l185;
  wire                when_SuperResolutionPart2_l195;
  wire                passPixels_fire_3;
  wire                when_SuperResolutionPart2_l200;
  wire                when_SuperResolutionPart2_l201;
  wire                passPixels_fire_4;
  wire                when_SuperResolutionPart2_l207;
  wire                when_SuperResolutionPart2_l208;
  wire                when_SuperResolutionPart2_l212;
  wire                controlStream_fire;
  wire                when_SuperResolutionPart2_l218;
  wire                when_SuperResolutionPart2_l220;
  wire                passPixels_fire_5;
  wire                when_SuperResolutionPart2_l224;
  wire                pixelsOut_fire;
  wire                when_SuperResolutionPart2_l234;
  wire                pixelsOut_fire_1;
  wire                when_SuperResolutionPart2_l235;
  wire                pixelsOut_fire_2;
  wire                pixelsOut_fire_3;
  wire                when_SuperResolutionPart2_l246;
  wire                passPixels_fire_6;
  wire                passPixels_fire_7;
  wire                passPixels_fire_8;
  wire                passPixels_fire_9;
  wire                passPixels_fire_10;
  wire                controlStream_fire_1;
  wire                pushing;
  wire                passPixels_fire_11;
  wire                controlStream_fire_2;
  wire                poping;
  wire                passPixels_fire_12;
  wire                controlStream_fire_3;
  wire                pushAndPoping;
  wire                mainAddrOneStream_s2mPipe_valid;
  reg                 mainAddrOneStream_s2mPipe_ready;
  wire       [10:0]   mainAddrOneStream_s2mPipe_payload;
  reg                 mainAddrOneStream_rValid;
  reg        [10:0]   mainAddrOneStream_rData;
  wire                mainAddrOneStream_s2mPipe_m2sPipe_valid;
  wire                mainAddrOneStream_s2mPipe_m2sPipe_ready;
  wire       [10:0]   mainAddrOneStream_s2mPipe_m2sPipe_payload;
  reg                 mainAddrOneStream_s2mPipe_rValid;
  reg        [10:0]   mainAddrOneStream_s2mPipe_rData;
  wire                when_Stream_l368_1;
  wire                CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_mainOnePixelStream_payload;
  reg                 CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_1;
  reg                 CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_mainOnePixelStream_payload_1;
  wire                readStage_mainOnePixelStream_valid;
  wire                readStage_mainOnePixelStream_ready;
  wire       [7:0]    readStage_mainOnePixelStream_payload;
  reg                 CICC1851_readStage_mainOnePixelStream_valid;
  reg        [7:0]    CICC1851_readStage_mainOnePixelStream_payload_2;
  wire                when_Stream_l368_2;
  wire                counterAddrOneStream_s2mPipe_valid;
  reg                 counterAddrOneStream_s2mPipe_ready;
  wire       [10:0]   counterAddrOneStream_s2mPipe_payload;
  reg                 counterAddrOneStream_rValid;
  reg        [10:0]   counterAddrOneStream_rData;
  wire                counterAddrOneStream_s2mPipe_m2sPipe_valid;
  wire                counterAddrOneStream_s2mPipe_m2sPipe_ready;
  wire       [10:0]   counterAddrOneStream_s2mPipe_m2sPipe_payload;
  reg                 counterAddrOneStream_s2mPipe_rValid;
  reg        [10:0]   counterAddrOneStream_s2mPipe_rData;
  wire                when_Stream_l368_3;
  wire                CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_counterOnePixelStream_payload;
  reg                 CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_2;
  reg                 CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_counterOnePixelStream_payload_1;
  wire                readStage_counterOnePixelStream_valid;
  wire                readStage_counterOnePixelStream_ready;
  wire       [7:0]    readStage_counterOnePixelStream_payload;
  reg                 CICC1851_readStage_counterOnePixelStream_valid;
  reg        [7:0]    CICC1851_readStage_counterOnePixelStream_payload_2;
  wire                when_Stream_l368_4;
  wire                mainAddrTwoStream_s2mPipe_valid;
  reg                 mainAddrTwoStream_s2mPipe_ready;
  wire       [10:0]   mainAddrTwoStream_s2mPipe_payload;
  reg                 mainAddrTwoStream_rValid;
  reg        [10:0]   mainAddrTwoStream_rData;
  wire                mainAddrTwoStream_s2mPipe_m2sPipe_valid;
  wire                mainAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire       [10:0]   mainAddrTwoStream_s2mPipe_m2sPipe_payload;
  reg                 mainAddrTwoStream_s2mPipe_rValid;
  reg        [10:0]   mainAddrTwoStream_s2mPipe_rData;
  wire                when_Stream_l368_5;
  wire                CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_mainTwoPixelStream_payload;
  reg                 CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_3;
  reg                 CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_mainTwoPixelStream_payload_1;
  wire                readStage_mainTwoPixelStream_valid;
  wire                readStage_mainTwoPixelStream_ready;
  wire       [7:0]    readStage_mainTwoPixelStream_payload;
  reg                 CICC1851_readStage_mainTwoPixelStream_valid;
  reg        [7:0]    CICC1851_readStage_mainTwoPixelStream_payload_2;
  wire                when_Stream_l368_6;
  wire                counterAddrTwoStream_s2mPipe_valid;
  reg                 counterAddrTwoStream_s2mPipe_ready;
  wire       [10:0]   counterAddrTwoStream_s2mPipe_payload;
  reg                 counterAddrTwoStream_rValid;
  reg        [10:0]   counterAddrTwoStream_rData;
  wire                counterAddrTwoStream_s2mPipe_m2sPipe_valid;
  wire                counterAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire       [10:0]   counterAddrTwoStream_s2mPipe_m2sPipe_payload;
  reg                 counterAddrTwoStream_s2mPipe_rValid;
  reg        [10:0]   counterAddrTwoStream_s2mPipe_rData;
  wire                when_Stream_l368_7;
  wire                CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_counterTwoPixelStream_payload;
  reg                 CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_4;
  reg                 CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_counterTwoPixelStream_payload_1;
  wire                readStage_counterTwoPixelStream_valid;
  wire                readStage_counterTwoPixelStream_ready;
  wire       [7:0]    readStage_counterTwoPixelStream_payload;
  reg                 CICC1851_readStage_counterTwoPixelStream_valid;
  reg        [7:0]    CICC1851_readStage_counterTwoPixelStream_payload_2;
  wire                when_Stream_l368_8;
  wire                oddAddrStream_s2mPipe_valid;
  reg                 oddAddrStream_s2mPipe_ready;
  wire       [10:0]   oddAddrStream_s2mPipe_payload;
  reg                 oddAddrStream_rValid;
  reg        [10:0]   oddAddrStream_rData;
  wire                oddAddrStream_s2mPipe_m2sPipe_valid;
  wire                oddAddrStream_s2mPipe_m2sPipe_ready;
  wire       [10:0]   oddAddrStream_s2mPipe_m2sPipe_payload;
  reg                 oddAddrStream_s2mPipe_rValid;
  reg        [10:0]   oddAddrStream_s2mPipe_rData;
  wire                when_Stream_l368_9;
  wire                CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_oddRowPixelStream_payload;
  reg                 CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_5;
  reg                 CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_oddRowPixelStream_payload_1;
  wire                readStage_oddRowPixelStream_valid;
  wire                readStage_oddRowPixelStream_ready;
  wire       [7:0]    readStage_oddRowPixelStream_payload;
  reg                 CICC1851_readStage_oddRowPixelStream_valid;
  reg        [7:0]    CICC1851_readStage_oddRowPixelStream_payload_2;
  wire                when_Stream_l368_10;
  wire                controlStream_s2mPipe_valid;
  reg                 controlStream_s2mPipe_ready;
  wire                controlStream_s2mPipe_payload_frameStart;
  wire                controlStream_s2mPipe_payload_rowEnd;
  wire                controlStream_s2mPipe_payload_passMode;
  wire                controlStream_s2mPipe_payload_passValid;
  wire       [2:0]    controlStream_s2mPipe_payload_onceMode;
  wire                controlStream_s2mPipe_payload_onceValid;
  wire                controlStream_s2mPipe_payload_mainCompare;
  wire                controlStream_s2mPipe_payload_counterCompare;
  wire       [7:0]    controlStream_s2mPipe_payload_mainDiff;
  wire       [7:0]    controlStream_s2mPipe_payload_counterDiff;
  wire                controlStream_s2mPipe_payload_twiceCompValid;
  wire       [2:0]    controlStream_s2mPipe_payload_twiceMode;
  wire                controlStream_s2mPipe_payload_inpValidFlag;
  wire                controlStream_s2mPipe_payload_oddValid;
  reg                 controlStream_rValid;
  reg                 controlStream_rData_frameStart;
  reg                 controlStream_rData_rowEnd;
  reg                 controlStream_rData_passMode;
  reg                 controlStream_rData_passValid;
  reg        [2:0]    controlStream_rData_onceMode;
  reg                 controlStream_rData_onceValid;
  reg                 controlStream_rData_mainCompare;
  reg                 controlStream_rData_counterCompare;
  reg        [7:0]    controlStream_rData_mainDiff;
  reg        [7:0]    controlStream_rData_counterDiff;
  reg                 controlStream_rData_twiceCompValid;
  reg        [2:0]    controlStream_rData_twiceMode;
  reg                 controlStream_rData_inpValidFlag;
  reg                 controlStream_rData_oddValid;
  wire                controlStream_s2mPipe_m2sPipe_valid;
  reg                 controlStream_s2mPipe_m2sPipe_ready;
  wire                controlStream_s2mPipe_m2sPipe_payload_frameStart;
  wire                controlStream_s2mPipe_m2sPipe_payload_rowEnd;
  wire                controlStream_s2mPipe_m2sPipe_payload_passMode;
  wire                controlStream_s2mPipe_m2sPipe_payload_passValid;
  wire       [2:0]    controlStream_s2mPipe_m2sPipe_payload_onceMode;
  wire                controlStream_s2mPipe_m2sPipe_payload_onceValid;
  wire                controlStream_s2mPipe_m2sPipe_payload_mainCompare;
  wire                controlStream_s2mPipe_m2sPipe_payload_counterCompare;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_payload_mainDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_payload_counterDiff;
  wire                controlStream_s2mPipe_m2sPipe_payload_twiceCompValid;
  wire       [2:0]    controlStream_s2mPipe_m2sPipe_payload_twiceMode;
  wire                controlStream_s2mPipe_m2sPipe_payload_inpValidFlag;
  wire                controlStream_s2mPipe_m2sPipe_payload_oddValid;
  reg                 controlStream_s2mPipe_rValid;
  reg                 controlStream_s2mPipe_rData_frameStart;
  reg                 controlStream_s2mPipe_rData_rowEnd;
  reg                 controlStream_s2mPipe_rData_passMode;
  reg                 controlStream_s2mPipe_rData_passValid;
  reg        [2:0]    controlStream_s2mPipe_rData_onceMode;
  reg                 controlStream_s2mPipe_rData_onceValid;
  reg                 controlStream_s2mPipe_rData_mainCompare;
  reg                 controlStream_s2mPipe_rData_counterCompare;
  reg        [7:0]    controlStream_s2mPipe_rData_mainDiff;
  reg        [7:0]    controlStream_s2mPipe_rData_counterDiff;
  reg                 controlStream_s2mPipe_rData_twiceCompValid;
  reg        [2:0]    controlStream_s2mPipe_rData_twiceMode;
  reg                 controlStream_s2mPipe_rData_inpValidFlag;
  reg                 controlStream_s2mPipe_rData_oddValid;
  wire                when_Stream_l368_11;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_valid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_ready;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_frameStart;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_rowEnd;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passMode;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passValid;
  wire       [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceMode;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceValid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainCompare;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterCompare;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDiff;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceCompValid;
  wire       [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceMode;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_inpValidFlag;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_oddValid;
  reg                 controlStream_s2mPipe_m2sPipe_rValid;
  reg                 controlStream_s2mPipe_m2sPipe_rData_frameStart;
  reg                 controlStream_s2mPipe_m2sPipe_rData_rowEnd;
  reg                 controlStream_s2mPipe_m2sPipe_rData_passMode;
  reg                 controlStream_s2mPipe_m2sPipe_rData_passValid;
  reg        [2:0]    controlStream_s2mPipe_m2sPipe_rData_onceMode;
  reg                 controlStream_s2mPipe_m2sPipe_rData_onceValid;
  reg                 controlStream_s2mPipe_m2sPipe_rData_mainCompare;
  reg                 controlStream_s2mPipe_m2sPipe_rData_counterCompare;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_rData_mainDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_rData_counterDiff;
  reg                 controlStream_s2mPipe_m2sPipe_rData_twiceCompValid;
  reg        [2:0]    controlStream_s2mPipe_m2sPipe_rData_twiceMode;
  reg                 controlStream_s2mPipe_m2sPipe_rData_inpValidFlag;
  reg                 controlStream_s2mPipe_m2sPipe_rData_oddValid;
  wire                when_Stream_l368_12;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_valid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_frameStart;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_rowEnd;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_passMode;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_passValid;
  wire       [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_onceMode;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_onceValid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainCompare;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterCompare;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterDiff;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_twiceCompValid;
  wire       [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_twiceMode;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_inpValidFlag;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_oddValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_frameStart;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_rowEnd;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_passMode;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_passValid;
  reg        [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_onceMode;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_onceValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainCompare;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterCompare;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterDiff;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_twiceCompValid;
  reg        [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_twiceMode;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_inpValidFlag;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_oddValid;
  wire                readStage_controlPipe_valid;
  wire                readStage_controlPipe_ready;
  wire                readStage_controlPipe_payload_frameStart;
  wire                readStage_controlPipe_payload_rowEnd;
  wire                readStage_controlPipe_payload_passMode;
  wire                readStage_controlPipe_payload_passValid;
  wire       [2:0]    readStage_controlPipe_payload_onceMode;
  wire                readStage_controlPipe_payload_onceValid;
  wire                readStage_controlPipe_payload_mainCompare;
  wire                readStage_controlPipe_payload_counterCompare;
  wire       [7:0]    readStage_controlPipe_payload_mainDiff;
  wire       [7:0]    readStage_controlPipe_payload_counterDiff;
  wire                readStage_controlPipe_payload_twiceCompValid;
  wire       [2:0]    readStage_controlPipe_payload_twiceMode;
  wire                readStage_controlPipe_payload_inpValidFlag;
  wire                readStage_controlPipe_payload_oddValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_frameStart;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_rowEnd;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_passMode;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_passValid;
  reg        [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_onceMode;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_onceValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainCompare;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterCompare;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterDiff;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_twiceCompValid;
  reg        [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_twiceMode;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_inpValidFlag;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_oddValid;
  wire                when_Stream_l368_13;
  wire                readStage_mainOnePixelStream_s2mPipe_valid;
  reg                 readStage_mainOnePixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_mainOnePixelStream_s2mPipe_payload;
  reg                 readStage_mainOnePixelStream_rValid;
  reg        [7:0]    readStage_mainOnePixelStream_rData;
  wire                compareStage_mainOnePixelStream_valid;
  wire                compareStage_mainOnePixelStream_ready;
  wire       [7:0]    compareStage_mainOnePixelStream_payload;
  reg                 readStage_mainOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_mainOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_14;
  wire                readStage_counterOnePixelStream_s2mPipe_valid;
  reg                 readStage_counterOnePixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_counterOnePixelStream_s2mPipe_payload;
  reg                 readStage_counterOnePixelStream_rValid;
  reg        [7:0]    readStage_counterOnePixelStream_rData;
  wire                compareStage_counterOnePixelStream_valid;
  wire                compareStage_counterOnePixelStream_ready;
  wire       [7:0]    compareStage_counterOnePixelStream_payload;
  reg                 readStage_counterOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_counterOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_15;
  wire                readStage_mainTwoPixelStream_s2mPipe_valid;
  reg                 readStage_mainTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_mainTwoPixelStream_s2mPipe_payload;
  reg                 readStage_mainTwoPixelStream_rValid;
  reg        [7:0]    readStage_mainTwoPixelStream_rData;
  wire                compareStage_mainTwoPixelStream_valid;
  wire                compareStage_mainTwoPixelStream_ready;
  wire       [7:0]    compareStage_mainTwoPixelStream_payload;
  reg                 readStage_mainTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_mainTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_16;
  wire                readStage_counterTwoPixelStream_s2mPipe_valid;
  reg                 readStage_counterTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_counterTwoPixelStream_s2mPipe_payload;
  reg                 readStage_counterTwoPixelStream_rValid;
  reg        [7:0]    readStage_counterTwoPixelStream_rData;
  wire                compareStage_counterTwoPixelStream_valid;
  wire                compareStage_counterTwoPixelStream_ready;
  wire       [7:0]    compareStage_counterTwoPixelStream_payload;
  reg                 readStage_counterTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_counterTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_17;
  wire                readStage_oddRowPixelStream_s2mPipe_valid;
  reg                 readStage_oddRowPixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_oddRowPixelStream_s2mPipe_payload;
  reg                 readStage_oddRowPixelStream_rValid;
  reg        [7:0]    readStage_oddRowPixelStream_rData;
  wire                compareStage_oddRowPixelStream_valid;
  wire                compareStage_oddRowPixelStream_ready;
  wire       [7:0]    compareStage_oddRowPixelStream_payload;
  reg                 readStage_oddRowPixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_oddRowPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_18;
  reg                 CICC1851_readStage_controlPipe_translated_payload_mainCompare;
  reg                 CICC1851_readStage_controlPipe_translated_payload_counterCompare;
  wire                when_SuperResolutionPart2_l290;
  wire                when_SuperResolutionPart2_l294;
  wire                when_SuperResolutionPart2_l298;
  wire                when_SuperResolutionPart2_l302;
  wire                when_SuperResolutionPart2_l313;
  wire                when_SuperResolutionPart2_l315;
  wire                when_SuperResolutionPart2_l319;
  wire                when_SuperResolutionPart2_l321;
  wire                when_SuperResolutionPart2_l326;
  wire                when_SuperResolutionPart2_l331;
  wire                readStage_controlPipe_translated_valid;
  wire                readStage_controlPipe_translated_ready;
  wire                readStage_controlPipe_translated_payload_frameStart;
  wire                readStage_controlPipe_translated_payload_rowEnd;
  wire                readStage_controlPipe_translated_payload_passMode;
  wire                readStage_controlPipe_translated_payload_passValid;
  wire       [2:0]    readStage_controlPipe_translated_payload_onceMode;
  wire                readStage_controlPipe_translated_payload_onceValid;
  wire                readStage_controlPipe_translated_payload_mainCompare;
  wire                readStage_controlPipe_translated_payload_counterCompare;
  wire       [7:0]    readStage_controlPipe_translated_payload_mainDiff;
  wire       [7:0]    readStage_controlPipe_translated_payload_counterDiff;
  wire                readStage_controlPipe_translated_payload_twiceCompValid;
  wire       [2:0]    readStage_controlPipe_translated_payload_twiceMode;
  wire                readStage_controlPipe_translated_payload_inpValidFlag;
  wire                readStage_controlPipe_translated_payload_oddValid;
  wire                readStage_controlPipe_translated_s2mPipe_valid;
  reg                 readStage_controlPipe_translated_s2mPipe_ready;
  wire                readStage_controlPipe_translated_s2mPipe_payload_frameStart;
  wire                readStage_controlPipe_translated_s2mPipe_payload_rowEnd;
  wire                readStage_controlPipe_translated_s2mPipe_payload_passMode;
  wire                readStage_controlPipe_translated_s2mPipe_payload_passValid;
  wire       [2:0]    readStage_controlPipe_translated_s2mPipe_payload_onceMode;
  wire                readStage_controlPipe_translated_s2mPipe_payload_onceValid;
  wire                readStage_controlPipe_translated_s2mPipe_payload_mainCompare;
  wire                readStage_controlPipe_translated_s2mPipe_payload_counterCompare;
  wire       [7:0]    readStage_controlPipe_translated_s2mPipe_payload_mainDiff;
  wire       [7:0]    readStage_controlPipe_translated_s2mPipe_payload_counterDiff;
  wire                readStage_controlPipe_translated_s2mPipe_payload_twiceCompValid;
  wire       [2:0]    readStage_controlPipe_translated_s2mPipe_payload_twiceMode;
  wire                readStage_controlPipe_translated_s2mPipe_payload_inpValidFlag;
  wire                readStage_controlPipe_translated_s2mPipe_payload_oddValid;
  reg                 readStage_controlPipe_translated_rValid;
  reg                 readStage_controlPipe_translated_rData_frameStart;
  reg                 readStage_controlPipe_translated_rData_rowEnd;
  reg                 readStage_controlPipe_translated_rData_passMode;
  reg                 readStage_controlPipe_translated_rData_passValid;
  reg        [2:0]    readStage_controlPipe_translated_rData_onceMode;
  reg                 readStage_controlPipe_translated_rData_onceValid;
  reg                 readStage_controlPipe_translated_rData_mainCompare;
  reg                 readStage_controlPipe_translated_rData_counterCompare;
  reg        [7:0]    readStage_controlPipe_translated_rData_mainDiff;
  reg        [7:0]    readStage_controlPipe_translated_rData_counterDiff;
  reg                 readStage_controlPipe_translated_rData_twiceCompValid;
  reg        [2:0]    readStage_controlPipe_translated_rData_twiceMode;
  reg                 readStage_controlPipe_translated_rData_inpValidFlag;
  reg                 readStage_controlPipe_translated_rData_oddValid;
  wire                compareStage_controlPipe_valid;
  wire                compareStage_controlPipe_ready;
  wire                compareStage_controlPipe_payload_frameStart;
  wire                compareStage_controlPipe_payload_rowEnd;
  wire                compareStage_controlPipe_payload_passMode;
  wire                compareStage_controlPipe_payload_passValid;
  wire       [2:0]    compareStage_controlPipe_payload_onceMode;
  wire                compareStage_controlPipe_payload_onceValid;
  wire                compareStage_controlPipe_payload_mainCompare;
  wire                compareStage_controlPipe_payload_counterCompare;
  wire       [7:0]    compareStage_controlPipe_payload_mainDiff;
  wire       [7:0]    compareStage_controlPipe_payload_counterDiff;
  wire                compareStage_controlPipe_payload_twiceCompValid;
  wire       [2:0]    compareStage_controlPipe_payload_twiceMode;
  wire                compareStage_controlPipe_payload_inpValidFlag;
  wire                compareStage_controlPipe_payload_oddValid;
  reg                 readStage_controlPipe_translated_s2mPipe_rValid;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_frameStart;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_rowEnd;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_passMode;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_passValid;
  reg        [2:0]    readStage_controlPipe_translated_s2mPipe_rData_onceMode;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_onceValid;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_mainCompare;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_counterCompare;
  reg        [7:0]    readStage_controlPipe_translated_s2mPipe_rData_mainDiff;
  reg        [7:0]    readStage_controlPipe_translated_s2mPipe_rData_counterDiff;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_twiceCompValid;
  reg        [2:0]    readStage_controlPipe_translated_s2mPipe_rData_twiceMode;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_inpValidFlag;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_oddValid;
  wire                when_Stream_l368_19;
  wire                compareStage_mainOnePixelStream_s2mPipe_valid;
  reg                 compareStage_mainOnePixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_mainOnePixelStream_s2mPipe_payload;
  reg                 compareStage_mainOnePixelStream_rValid;
  reg        [7:0]    compareStage_mainOnePixelStream_rData;
  wire                diffStage_mainOnePixelStream_valid;
  wire                diffStage_mainOnePixelStream_ready;
  wire       [7:0]    diffStage_mainOnePixelStream_payload;
  reg                 compareStage_mainOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_mainOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_20;
  wire                compareStage_counterOnePixelStream_s2mPipe_valid;
  reg                 compareStage_counterOnePixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_counterOnePixelStream_s2mPipe_payload;
  reg                 compareStage_counterOnePixelStream_rValid;
  reg        [7:0]    compareStage_counterOnePixelStream_rData;
  wire                diffStage_counterOnePixelStream_valid;
  wire                diffStage_counterOnePixelStream_ready;
  wire       [7:0]    diffStage_counterOnePixelStream_payload;
  reg                 compareStage_counterOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_counterOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_21;
  wire                compareStage_mainTwoPixelStream_s2mPipe_valid;
  reg                 compareStage_mainTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_mainTwoPixelStream_s2mPipe_payload;
  reg                 compareStage_mainTwoPixelStream_rValid;
  reg        [7:0]    compareStage_mainTwoPixelStream_rData;
  wire                diffStage_mainTwoPixelStream_valid;
  wire                diffStage_mainTwoPixelStream_ready;
  wire       [7:0]    diffStage_mainTwoPixelStream_payload;
  reg                 compareStage_mainTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_mainTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_22;
  wire                compareStage_counterTwoPixelStream_s2mPipe_valid;
  reg                 compareStage_counterTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_counterTwoPixelStream_s2mPipe_payload;
  reg                 compareStage_counterTwoPixelStream_rValid;
  reg        [7:0]    compareStage_counterTwoPixelStream_rData;
  wire                diffStage_counterTwoPixelStream_valid;
  wire                diffStage_counterTwoPixelStream_ready;
  wire       [7:0]    diffStage_counterTwoPixelStream_payload;
  reg                 compareStage_counterTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_counterTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_23;
  wire                compareStage_oddRowPixelStream_s2mPipe_valid;
  reg                 compareStage_oddRowPixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_oddRowPixelStream_s2mPipe_payload;
  reg                 compareStage_oddRowPixelStream_rValid;
  reg        [7:0]    compareStage_oddRowPixelStream_rData;
  wire                diffStage_oddRowPixelStream_valid;
  wire                diffStage_oddRowPixelStream_ready;
  wire       [7:0]    diffStage_oddRowPixelStream_payload;
  reg                 compareStage_oddRowPixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_oddRowPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_24;
  reg        [7:0]    CICC1851_compareStage_controlPipe_translated_payload_mainDiff;
  reg        [7:0]    CICC1851_compareStage_controlPipe_translated_payload_counterDiff;
  wire                compareStage_controlPipe_translated_valid;
  wire                compareStage_controlPipe_translated_ready;
  wire                compareStage_controlPipe_translated_payload_frameStart;
  wire                compareStage_controlPipe_translated_payload_rowEnd;
  wire                compareStage_controlPipe_translated_payload_passMode;
  wire                compareStage_controlPipe_translated_payload_passValid;
  wire       [2:0]    compareStage_controlPipe_translated_payload_onceMode;
  wire                compareStage_controlPipe_translated_payload_onceValid;
  wire                compareStage_controlPipe_translated_payload_mainCompare;
  wire                compareStage_controlPipe_translated_payload_counterCompare;
  wire       [7:0]    compareStage_controlPipe_translated_payload_mainDiff;
  wire       [7:0]    compareStage_controlPipe_translated_payload_counterDiff;
  wire                compareStage_controlPipe_translated_payload_twiceCompValid;
  wire       [2:0]    compareStage_controlPipe_translated_payload_twiceMode;
  wire                compareStage_controlPipe_translated_payload_inpValidFlag;
  wire                compareStage_controlPipe_translated_payload_oddValid;
  wire                compareStage_controlPipe_translated_s2mPipe_valid;
  reg                 compareStage_controlPipe_translated_s2mPipe_ready;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_frameStart;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_rowEnd;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_passMode;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_passValid;
  wire       [2:0]    compareStage_controlPipe_translated_s2mPipe_payload_onceMode;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_onceValid;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_mainCompare;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_counterCompare;
  wire       [7:0]    compareStage_controlPipe_translated_s2mPipe_payload_mainDiff;
  wire       [7:0]    compareStage_controlPipe_translated_s2mPipe_payload_counterDiff;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_twiceCompValid;
  wire       [2:0]    compareStage_controlPipe_translated_s2mPipe_payload_twiceMode;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_inpValidFlag;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_oddValid;
  reg                 compareStage_controlPipe_translated_rValid;
  reg                 compareStage_controlPipe_translated_rData_frameStart;
  reg                 compareStage_controlPipe_translated_rData_rowEnd;
  reg                 compareStage_controlPipe_translated_rData_passMode;
  reg                 compareStage_controlPipe_translated_rData_passValid;
  reg        [2:0]    compareStage_controlPipe_translated_rData_onceMode;
  reg                 compareStage_controlPipe_translated_rData_onceValid;
  reg                 compareStage_controlPipe_translated_rData_mainCompare;
  reg                 compareStage_controlPipe_translated_rData_counterCompare;
  reg        [7:0]    compareStage_controlPipe_translated_rData_mainDiff;
  reg        [7:0]    compareStage_controlPipe_translated_rData_counterDiff;
  reg                 compareStage_controlPipe_translated_rData_twiceCompValid;
  reg        [2:0]    compareStage_controlPipe_translated_rData_twiceMode;
  reg                 compareStage_controlPipe_translated_rData_inpValidFlag;
  reg                 compareStage_controlPipe_translated_rData_oddValid;
  wire                diffStage_controlPipe_valid;
  wire                diffStage_controlPipe_ready;
  wire                diffStage_controlPipe_payload_frameStart;
  wire                diffStage_controlPipe_payload_rowEnd;
  wire                diffStage_controlPipe_payload_passMode;
  wire                diffStage_controlPipe_payload_passValid;
  wire       [2:0]    diffStage_controlPipe_payload_onceMode;
  wire                diffStage_controlPipe_payload_onceValid;
  wire                diffStage_controlPipe_payload_mainCompare;
  wire                diffStage_controlPipe_payload_counterCompare;
  wire       [7:0]    diffStage_controlPipe_payload_mainDiff;
  wire       [7:0]    diffStage_controlPipe_payload_counterDiff;
  wire                diffStage_controlPipe_payload_twiceCompValid;
  wire       [2:0]    diffStage_controlPipe_payload_twiceMode;
  wire                diffStage_controlPipe_payload_inpValidFlag;
  wire                diffStage_controlPipe_payload_oddValid;
  reg                 compareStage_controlPipe_translated_s2mPipe_rValid;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_frameStart;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_rowEnd;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_passMode;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_passValid;
  reg        [2:0]    compareStage_controlPipe_translated_s2mPipe_rData_onceMode;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_onceValid;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_mainCompare;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_counterCompare;
  reg        [7:0]    compareStage_controlPipe_translated_s2mPipe_rData_mainDiff;
  reg        [7:0]    compareStage_controlPipe_translated_s2mPipe_rData_counterDiff;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_twiceCompValid;
  reg        [2:0]    compareStage_controlPipe_translated_s2mPipe_rData_twiceMode;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_inpValidFlag;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_oddValid;
  wire                when_Stream_l368_25;
  wire                diffStage_mainOnePixelStream_s2mPipe_valid;
  reg                 diffStage_mainOnePixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_mainOnePixelStream_s2mPipe_payload;
  reg                 diffStage_mainOnePixelStream_rValid;
  reg        [7:0]    diffStage_mainOnePixelStream_rData;
  wire                resultStage_mainOnePixelStream_valid;
  wire                resultStage_mainOnePixelStream_ready;
  wire       [7:0]    resultStage_mainOnePixelStream_payload;
  reg                 diffStage_mainOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_mainOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_26;
  wire                diffStage_counterOnePixelStream_s2mPipe_valid;
  reg                 diffStage_counterOnePixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_counterOnePixelStream_s2mPipe_payload;
  reg                 diffStage_counterOnePixelStream_rValid;
  reg        [7:0]    diffStage_counterOnePixelStream_rData;
  wire                resultStage_counterOnePixelStream_valid;
  wire                resultStage_counterOnePixelStream_ready;
  wire       [7:0]    resultStage_counterOnePixelStream_payload;
  reg                 diffStage_counterOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_counterOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_27;
  wire                diffStage_mainTwoPixelStream_s2mPipe_valid;
  reg                 diffStage_mainTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_mainTwoPixelStream_s2mPipe_payload;
  reg                 diffStage_mainTwoPixelStream_rValid;
  reg        [7:0]    diffStage_mainTwoPixelStream_rData;
  wire                resultStage_mainTwoPixelStream_valid;
  wire                resultStage_mainTwoPixelStream_ready;
  wire       [7:0]    resultStage_mainTwoPixelStream_payload;
  reg                 diffStage_mainTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_mainTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_28;
  wire                diffStage_counterTwoPixelStream_s2mPipe_valid;
  reg                 diffStage_counterTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_counterTwoPixelStream_s2mPipe_payload;
  reg                 diffStage_counterTwoPixelStream_rValid;
  reg        [7:0]    diffStage_counterTwoPixelStream_rData;
  wire                resultStage_counterTwoPixelStream_valid;
  wire                resultStage_counterTwoPixelStream_ready;
  wire       [7:0]    resultStage_counterTwoPixelStream_payload;
  reg                 diffStage_counterTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_counterTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_29;
  wire                diffStage_oddRowPixelStream_s2mPipe_valid;
  reg                 diffStage_oddRowPixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_oddRowPixelStream_s2mPipe_payload;
  reg                 diffStage_oddRowPixelStream_rValid;
  reg        [7:0]    diffStage_oddRowPixelStream_rData;
  wire                resultStage_oddRowPixelStream_valid;
  wire                resultStage_oddRowPixelStream_ready;
  wire       [7:0]    resultStage_oddRowPixelStream_payload;
  reg                 diffStage_oddRowPixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_oddRowPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_30;
  wire       [2:0]    CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceMode;
  wire                CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceValid;
  wire       [7:0]    CICC1851_when_SuperResolutionPart2_l419;
  wire       [7:0]    CICC1851_when_SuperResolutionPart2_l428;
  wire                CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceCompValid;
  wire       [2:0]    CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceMode;
  reg                 CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag;
  wire                when_SuperResolutionPart2_l419;
  wire                when_SuperResolutionPart2_l420;
  wire                when_SuperResolutionPart2_l421;
  wire                when_SuperResolutionPart2_l422;
  wire                when_SuperResolutionPart2_l428;
  wire                when_SuperResolutionPart2_l429;
  wire                when_SuperResolutionPart2_l430;
  wire                when_SuperResolutionPart2_l431;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_valid;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_ready;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_payload_frameStart;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_payload_rowEnd;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_payload_passMode;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_payload_passValid;
  wire       [2:0]    diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceMode;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceValid;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_payload_mainCompare;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_payload_counterCompare;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_translated_payload_mainDiff;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_translated_payload_counterDiff;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceCompValid;
  wire       [2:0]    diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceMode;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_payload_oddValid;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_valid;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_ready;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_frameStart;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_rowEnd;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_passMode;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_passValid;
  wire       [2:0]    diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_onceMode;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_onceValid;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_mainCompare;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_counterCompare;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_mainDiff;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_counterDiff;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_twiceCompValid;
  wire       [2:0]    diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_twiceMode;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_inpValidFlag;
  wire                diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_oddValid;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_rValid;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_rData_frameStart;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_rData_rowEnd;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_rData_passMode;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_rData_passValid;
  reg        [2:0]    diffStage_controlPipe_fork_io_outputs_0_translated_rData_onceMode;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_rData_onceValid;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_rData_mainCompare;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_rData_counterCompare;
  reg        [7:0]    diffStage_controlPipe_fork_io_outputs_0_translated_rData_mainDiff;
  reg        [7:0]    diffStage_controlPipe_fork_io_outputs_0_translated_rData_counterDiff;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_rData_twiceCompValid;
  reg        [2:0]    diffStage_controlPipe_fork_io_outputs_0_translated_rData_twiceMode;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_rData_inpValidFlag;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_rData_oddValid;
  wire                resultStage_controlPipe_valid;
  wire                resultStage_controlPipe_ready;
  wire                resultStage_controlPipe_payload_frameStart;
  wire                resultStage_controlPipe_payload_rowEnd;
  wire                resultStage_controlPipe_payload_passMode;
  wire                resultStage_controlPipe_payload_passValid;
  wire       [2:0]    resultStage_controlPipe_payload_onceMode;
  wire                resultStage_controlPipe_payload_onceValid;
  wire                resultStage_controlPipe_payload_mainCompare;
  wire                resultStage_controlPipe_payload_counterCompare;
  wire       [7:0]    resultStage_controlPipe_payload_mainDiff;
  wire       [7:0]    resultStage_controlPipe_payload_counterDiff;
  wire                resultStage_controlPipe_payload_twiceCompValid;
  wire       [2:0]    resultStage_controlPipe_payload_twiceMode;
  wire                resultStage_controlPipe_payload_inpValidFlag;
  wire                resultStage_controlPipe_payload_oddValid;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rValid;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_frameStart;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_rowEnd;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_passMode;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_passValid;
  reg        [2:0]    diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_onceMode;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_onceValid;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_mainCompare;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_counterCompare;
  reg        [7:0]    diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_mainDiff;
  reg        [7:0]    diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_counterDiff;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_twiceCompValid;
  reg        [2:0]    diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_twiceMode;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_inpValidFlag;
  reg                 diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_oddValid;
  wire                when_Stream_l368_31;
  wire                resultStage_pixelStream_valid;
  wire                resultStage_pixelStream_ready;
  reg        [7:0]    resultStage_pixelStream_payload;
  wire                when_SuperResolutionPart2_l451;
  wire                when_SuperResolutionPart2_l455;
  wire                when_SuperResolutionPart2_l459;
  wire                when_SuperResolutionPart2_l463;
  wire                when_SuperResolutionPart2_l474;
  wire                when_SuperResolutionPart2_l477;
  wire                when_SuperResolutionPart2_l482;
  wire                when_SuperResolutionPart2_l485;
  wire                when_SuperResolutionPart2_l491;
  wire                when_SuperResolutionPart2_l496;
  wire                resultStage_pixelStream_s2mPipe_valid;
  reg                 resultStage_pixelStream_s2mPipe_ready;
  wire       [7:0]    resultStage_pixelStream_s2mPipe_payload;
  reg                 resultStage_pixelStream_rValid;
  reg        [7:0]    resultStage_pixelStream_rData;
  wire                resultStage_resultStream_valid;
  wire                resultStage_resultStream_ready;
  wire       [7:0]    resultStage_resultStream_payload;
  reg                 resultStage_pixelStream_s2mPipe_rValid;
  reg        [7:0]    resultStage_pixelStream_s2mPipe_rData;
  wire                when_Stream_l368_32;
  wire                CICC1851_resultStage_mainOnePixelStream_ready;
  reg                 CICC1851_resultStage_mainOnePixelStream_ready_1;
  wire                CICC1851_resultStage_mainOnePixelStream_ready_2;
  wire                when_Stream_l438;
  reg                 resultsJoin_valid;
  wire                resultsJoin_ready;
  wire                pixelsStream_valid;
  wire                pixelsStream_ready;
  wire       [7:0]    pixelsStream_payload_pixel;
  wire                pixelsStream_payload_frameStart;
  wire                pixelsStream_payload_rowEnd;
  wire                pixelsStream_payload_inpValid;
  wire                pixelsStream_s2mPipe_valid;
  reg                 pixelsStream_s2mPipe_ready;
  wire       [7:0]    pixelsStream_s2mPipe_payload_pixel;
  wire                pixelsStream_s2mPipe_payload_frameStart;
  wire                pixelsStream_s2mPipe_payload_rowEnd;
  wire                pixelsStream_s2mPipe_payload_inpValid;
  reg                 pixelsStream_rValid;
  reg        [7:0]    pixelsStream_rData_pixel;
  reg                 pixelsStream_rData_frameStart;
  reg                 pixelsStream_rData_rowEnd;
  reg                 pixelsStream_rData_inpValid;
  wire                pixelsStream_s2mPipe_m2sPipe_valid;
  wire                pixelsStream_s2mPipe_m2sPipe_ready;
  wire       [7:0]    pixelsStream_s2mPipe_m2sPipe_payload_pixel;
  wire                pixelsStream_s2mPipe_m2sPipe_payload_frameStart;
  wire                pixelsStream_s2mPipe_m2sPipe_payload_rowEnd;
  wire                pixelsStream_s2mPipe_m2sPipe_payload_inpValid;
  reg                 pixelsStream_s2mPipe_rValid;
  reg        [7:0]    pixelsStream_s2mPipe_rData_pixel;
  reg                 pixelsStream_s2mPipe_rData_frameStart;
  reg                 pixelsStream_s2mPipe_rData_rowEnd;
  reg                 pixelsStream_s2mPipe_rData_inpValid;
  wire                when_Stream_l368_33;
  wire                controlStateMachine_wantExit;
  reg                 controlStateMachine_wantStart;
  wire                controlStateMachine_wantKill;
  wire                when_SuperResolutionPart2_l761;
  wire                controlStream_fire_4;
  wire                when_SuperResolutionPart2_l763;
  wire                controlStream_fire_5;
  wire                when_SuperResolutionPart2_l764;
  wire                controlStream_fire_6;
  wire                when_SuperResolutionPart2_l766;
  wire                controlStream_fire_7;
  wire                when_SuperResolutionPart2_l783;
  wire                when_SuperResolutionPart2_l785;
  wire                when_SuperResolutionPart2_l787;
  wire                when_SuperResolutionPart2_l789;
  wire                when_SuperResolutionPart2_l793;
  wire                when_SuperResolutionPart2_l796;
  wire                when_SuperResolutionPart2_l799;
  wire                when_SuperResolutionPart2_l802;
  reg        [2:0]    controlStateMachine_stateReg;
  reg        [2:0]    controlStateMachine_stateNext;
  wire                passPixels_fire_13;
  wire                passPixels_fire_14;
  wire                passPixels_fire_15;
  wire                passPixels_fire_16;
  wire                when_SuperResolutionPart2_l560;
  wire                controlStream_fire_8;
  wire                passPixels_fire_17;
  wire                when_SuperResolutionPart2_l573;
  wire                passPixels_fire_18;
  wire                when_SuperResolutionPart2_l578;
  wire                when_SuperResolutionPart2_l585;
  wire                when_SuperResolutionPart2_l588;
  wire                passPixels_fire_19;
  wire                when_SuperResolutionPart2_l590;
  wire                when_SuperResolutionPart2_l602;
  wire                when_SuperResolutionPart2_l603;
  wire                when_SuperResolutionPart2_l605;
  wire                when_SuperResolutionPart2_l606;
  wire                when_SuperResolutionPart2_l609;
  wire                controlStream_fire_9;
  wire                when_SuperResolutionPart2_l630;
  wire                controlStream_fire_10;
  wire                passPixels_fire_20;
  wire                when_SuperResolutionPart2_l642;
  wire                passPixels_fire_21;
  wire                when_SuperResolutionPart2_l647;
  wire                passPixels_fire_22;
  wire                when_SuperResolutionPart2_l653;
  wire                passPixels_fire_23;
  wire                when_SuperResolutionPart2_l662;
  wire                when_SuperResolutionPart2_l667;
  wire                when_SuperResolutionPart2_l668;
  wire                controlStream_fire_11;
  `ifndef SYNTHESIS
  reg [39:0] controlStateMachine_stateReg_string;
  reg [39:0] controlStateMachine_stateNext_string;
  `endif

  reg [7:0] lineBufferOne [0:1919];
  reg [7:0] lineBufferTwo [0:1919];
  reg [7:0] lineBufferOdd [0:1919];

  assign CICC1851_bufferRowCount_valueNext_1 = bufferRowCount_willIncrement;
  assign CICC1851_bufferRowCount_valueNext = {10'd0, CICC1851_bufferRowCount_valueNext_1};
  assign CICC1851_bufferWAddr_valueNext_1 = bufferWAddr_willIncrement;
  assign CICC1851_bufferWAddr_valueNext = {10'd0, CICC1851_bufferWAddr_valueNext_1};
  assign CICC1851_outPixelAddr_valueNext_1 = outPixelAddr_willIncrement;
  assign CICC1851_outPixelAddr_valueNext = {11'd0, CICC1851_outPixelAddr_valueNext_1};
  assign CICC1851_outRowCount_valueNext_1 = outRowCount_willIncrement;
  assign CICC1851_outRowCount_valueNext = {11'd0, CICC1851_outRowCount_valueNext_1};
  assign CICC1851_alreadySendRow_valueNext_1 = alreadySendRow_willIncrement;
  assign CICC1851_alreadySendRow_valueNext = {11'd0, CICC1851_alreadySendRow_valueNext_1};
  assign CICC1851_alreadySendCountInRow_valueNext_1 = alreadySendCountInRow_willIncrement;
  assign CICC1851_alreadySendCountInRow_valueNext = {11'd0, CICC1851_alreadySendCountInRow_valueNext_1};
  assign CICC1851_mainAddrOne = (outPixelAddr_value / 2'b10);
  assign CICC1851_counterAddrOne = (outPixelAddr_value / 2'b10);
  assign CICC1851_mainAddrTwo = (outPixelAddr_value / 2'b10);
  assign CICC1851_counterAddrTwo = (outPixelAddr_value / 2'b10);
  assign CICC1851_oddAddr = (outPixelAddr_value / 2'b10);
  assign CICC1851_when_SuperResolutionPart2_l181 = {1'd0, bufferWAddr_value};
  assign CICC1851_when_SuperResolutionPart2_l181_1 = (CICC1851_when_SuperResolutionPart2_l181_2 - 12'h002);
  assign CICC1851_when_SuperResolutionPart2_l181_2 = (2'b10 * bmpWidth);
  assign CICC1851_when_SuperResolutionPart2_l182 = {1'd0, bufferRowCount_value};
  assign CICC1851_when_SuperResolutionPart2_l182_1 = (CICC1851_when_SuperResolutionPart2_l182_2 - 12'h002);
  assign CICC1851_when_SuperResolutionPart2_l182_2 = (2'b10 * bmpHeight);
  assign CICC1851_when_SuperResolutionPart2_l195 = (bufferRowCount_value % 2'b10);
  assign CICC1851_when_SuperResolutionPart2_l218 = (outRowCount_value % 3'b100);
  assign CICC1851_when_SuperResolutionPart2_l234 = {1'd0, alreadySendCountInRow_value};
  assign CICC1851_when_SuperResolutionPart2_l234_1 = (CICC1851_when_SuperResolutionPart2_l234_2 - 13'h0002);
  assign CICC1851_when_SuperResolutionPart2_l234_2 = (3'b100 * bmpWidth);
  assign CICC1851_when_SuperResolutionPart2_l235 = {1'd0, alreadySendRow_value};
  assign CICC1851_when_SuperResolutionPart2_l235_1 = (CICC1851_when_SuperResolutionPart2_l235_2 - 13'h0002);
  assign CICC1851_when_SuperResolutionPart2_l235_2 = (3'b100 * bmpHeight);
  assign CICC1851_resultStage_pixelStream_payload = (CICC1851_resultStage_pixelStream_payload_1 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_1 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_2 = (CICC1851_resultStage_pixelStream_payload_3 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_3 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_4 = (CICC1851_resultStage_pixelStream_payload_5 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_5 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_mainTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_6 = (CICC1851_resultStage_pixelStream_payload_7 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_7 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_mainOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_8 = (CICC1851_resultStage_pixelStream_payload_9 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_9 = ({1'b0,diffStage_counterOnePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_10 = (CICC1851_resultStage_pixelStream_payload_11 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_11 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_mainTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_12 = (CICC1851_resultStage_pixelStream_payload_13 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_13 = ({1'b0,diffStage_counterOnePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_14 = (CICC1851_resultStage_pixelStream_payload_15 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_15 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_mainTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_16 = (CICC1851_resultStage_pixelStream_payload_17 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_17 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_18 = (CICC1851_resultStage_pixelStream_payload_19 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_19 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_when_SuperResolutionPart2_l763 = {1'd0, outPixelAddr_value};
  assign CICC1851_when_SuperResolutionPart2_l763_1 = (CICC1851_when_SuperResolutionPart2_l763_2 - 13'h0002);
  assign CICC1851_when_SuperResolutionPart2_l763_2 = (3'b100 * bmpWidth);
  assign CICC1851_when_SuperResolutionPart2_l764 = {1'd0, outRowCount_value};
  assign CICC1851_when_SuperResolutionPart2_l764_1 = (CICC1851_when_SuperResolutionPart2_l764_2 - 13'h0002);
  assign CICC1851_when_SuperResolutionPart2_l764_2 = (3'b100 * bmpHeight);
  assign CICC1851_when_SuperResolutionPart2_l783 = (outRowCount_value % 3'b100);
  assign CICC1851_when_SuperResolutionPart2_l785 = (outRowCount_value % 3'b100);
  assign CICC1851_when_SuperResolutionPart2_l787 = (outRowCount_value % 3'b100);
  assign CICC1851_when_SuperResolutionPart2_l789 = (outRowCount_value % 3'b100);
  assign CICC1851_when_SuperResolutionPart2_l793 = (outPixelAddr_value % 3'b100);
  assign CICC1851_when_SuperResolutionPart2_l796 = (outPixelAddr_value % 3'b100);
  assign CICC1851_when_SuperResolutionPart2_l799 = (outPixelAddr_value % 3'b100);
  assign CICC1851_when_SuperResolutionPart2_l802 = (outPixelAddr_value % 3'b100);
  assign CICC1851_when_SuperResolutionPart2_l560 = (2'b10 * bufferWAddr_value);
  assign CICC1851_when_SuperResolutionPart2_l560_1 = {1'd0, outPixelAddr_value};
  assign CICC1851_when_SuperResolutionPart2_l602 = (2'b10 * bufferWAddr_value);
  assign CICC1851_when_SuperResolutionPart2_l602_1 = (CICC1851_when_SuperResolutionPart2_l602_2 + {1'b0,outPixelAddr_value});
  assign CICC1851_when_SuperResolutionPart2_l602_3 = {1'b0,2'b10};
  assign CICC1851_when_SuperResolutionPart2_l602_2 = {10'd0, CICC1851_when_SuperResolutionPart2_l602_3};
  assign CICC1851_when_SuperResolutionPart2_l603 = (2'b10 * bufferWAddr_value);
  assign CICC1851_when_SuperResolutionPart2_l603_1 = {1'd0, outPixelAddr_value};
  assign CICC1851_when_SuperResolutionPart2_l605 = (2'b10 * bufferWAddr_value);
  assign CICC1851_when_SuperResolutionPart2_l605_1 = (CICC1851_when_SuperResolutionPart2_l605_2 + {1'b0,outPixelAddr_value});
  assign CICC1851_when_SuperResolutionPart2_l605_3 = {1'b0,2'b11};
  assign CICC1851_when_SuperResolutionPart2_l605_2 = {10'd0, CICC1851_when_SuperResolutionPart2_l605_3};
  assign CICC1851_when_SuperResolutionPart2_l606 = (2'b10 * bufferWAddr_value);
  assign CICC1851_when_SuperResolutionPart2_l606_1 = (CICC1851_when_SuperResolutionPart2_l606_2 + {1'b0,outPixelAddr_value});
  assign CICC1851_when_SuperResolutionPart2_l606_3 = {1'b0,1'b1};
  assign CICC1851_when_SuperResolutionPart2_l606_2 = {11'd0, CICC1851_when_SuperResolutionPart2_l606_3};
  assign CICC1851_when_SuperResolutionPart2_l609 = (outPixelAddr_value % 2'b10);
  assign CICC1851_mainAddrOne_1 = (CICC1851_mainAddrOne_2 / 2'b10);
  assign CICC1851_mainAddrOne_2 = (outPixelAddr_value - 12'h002);
  assign CICC1851_mainAddrTwo_1 = (CICC1851_mainAddrTwo_2 / 2'b10);
  assign CICC1851_mainAddrTwo_2 = (outPixelAddr_value - 12'h002);
  assign CICC1851_when_SuperResolutionPart2_l667 = (CICC1851_when_SuperResolutionPart2_l667_1 - 13'h0002);
  assign CICC1851_when_SuperResolutionPart2_l667_1 = (2'b10 * bufferWAddr_value);
  assign CICC1851_when_SuperResolutionPart2_l667_2 = (CICC1851_when_SuperResolutionPart2_l667_3 + {1'b0,outPixelAddr_value});
  assign CICC1851_when_SuperResolutionPart2_l667_4 = {1'b0,1'b1};
  assign CICC1851_when_SuperResolutionPart2_l667_3 = {11'd0, CICC1851_when_SuperResolutionPart2_l667_4};
  assign CICC1851_when_SuperResolutionPart2_l668 = (2'b10 * bufferWAddr_value);
  assign CICC1851_when_SuperResolutionPart2_l668_1 = (CICC1851_when_SuperResolutionPart2_l668_2 + {1'b0,outPixelAddr_value});
  assign CICC1851_when_SuperResolutionPart2_l668_3 = {1'b0,1'b1};
  assign CICC1851_when_SuperResolutionPart2_l668_2 = {11'd0, CICC1851_when_SuperResolutionPart2_l668_3};
  assign CICC1851_mainAddrOne_3 = (CICC1851_mainAddrOne_4 / 2'b10);
  assign CICC1851_mainAddrOne_4 = (outPixelAddr_value - 12'h002);
  assign CICC1851_mainAddrTwo_3 = (CICC1851_mainAddrTwo_4 / 2'b10);
  assign CICC1851_mainAddrTwo_4 = (outPixelAddr_value - 12'h002);
  assign CICC1851_controls_onceMode = 2'b10;
  assign CICC1851_controls_onceMode_1 = 2'b11;
  assign CICC1851_mainAddrOne_5 = (CICC1851_mainAddrOne_6 / 2'b10);
  assign CICC1851_mainAddrOne_6 = (outPixelAddr_value - 12'h003);
  assign CICC1851_counterAddrOne_1 = (CICC1851_counterAddrOne_2 / 2'b10);
  assign CICC1851_counterAddrOne_2 = (outPixelAddr_value - 12'h003);
  assign CICC1851_counterAddrOne_3 = (CICC1851_counterAddrOne_4 / 2'b10);
  assign CICC1851_counterAddrOne_4 = (12'h001 + outPixelAddr_value);
  assign CICC1851_controls_onceMode_2 = 1'b1;
  assign CICC1851_mainAddrTwo_5 = (CICC1851_mainAddrTwo_6 / 2'b10);
  assign CICC1851_mainAddrTwo_6 = (outPixelAddr_value - 12'h003);
  assign CICC1851_counterAddrTwo_1 = (CICC1851_counterAddrTwo_2 / 2'b10);
  assign CICC1851_counterAddrTwo_2 = (outPixelAddr_value - 12'h003);
  assign CICC1851_counterAddrTwo_3 = (CICC1851_counterAddrTwo_4 / 2'b10);
  assign CICC1851_counterAddrTwo_4 = (12'h001 + outPixelAddr_value);
  assign CICC1851_mainAddrOne_7 = (CICC1851_mainAddrOne_8 / 2'b10);
  assign CICC1851_mainAddrOne_8 = (outPixelAddr_value - 12'h003);
  assign CICC1851_mainAddrOne_9 = (CICC1851_mainAddrOne_10 / 2'b10);
  assign CICC1851_mainAddrOne_10 = (outPixelAddr_value - 12'h003);
  assign CICC1851_counterAddrOne_5 = (CICC1851_counterAddrOne_6 / 2'b10);
  assign CICC1851_counterAddrOne_6 = (CICC1851_counterAddrOne_7 + {1'b0,outPixelAddr_value});
  assign CICC1851_counterAddrOne_8 = {1'b0,1'b1};
  assign CICC1851_counterAddrOne_7 = {11'd0, CICC1851_counterAddrOne_8};
  assign CICC1851_controls_twiceMode = 2'b10;
  assign CICC1851_mainAddrTwo_7 = (CICC1851_mainAddrTwo_8 / 2'b10);
  assign CICC1851_mainAddrTwo_8 = (outPixelAddr_value - 12'h003);
  assign CICC1851_controls_twiceMode_1 = 2'b11;
  assign CICC1851_mainAddrTwo_9 = (CICC1851_mainAddrTwo_10 / 2'b10);
  assign CICC1851_mainAddrTwo_10 = (outPixelAddr_value - 12'h003);
  assign CICC1851_counterAddrTwo_5 = (CICC1851_counterAddrTwo_6 / 2'b10);
  assign CICC1851_counterAddrTwo_6 = (CICC1851_counterAddrTwo_7 + {1'b0,outPixelAddr_value});
  assign CICC1851_counterAddrTwo_8 = {1'b0,1'b1};
  assign CICC1851_counterAddrTwo_7 = {11'd0, CICC1851_counterAddrTwo_8};
  assign CICC1851_mainAddrOne_11 = (CICC1851_mainAddrOne_12 / 2'b10);
  assign CICC1851_mainAddrOne_12 = (outPixelAddr_value - 12'h003);
  assign CICC1851_counterAddrTwo_9 = (CICC1851_counterAddrTwo_10 / 2'b10);
  assign CICC1851_counterAddrTwo_10 = (outPixelAddr_value - 12'h003);
  assign CICC1851_mainAddrTwo_11 = (CICC1851_mainAddrTwo_12 / 2'b10);
  assign CICC1851_mainAddrTwo_12 = (outPixelAddr_value - 12'h003);
  assign CICC1851_counterAddrOne_9 = (CICC1851_counterAddrOne_10 / 2'b10);
  assign CICC1851_counterAddrOne_10 = (outPixelAddr_value - 12'h003);
  assign CICC1851_mainAddrTwo_13 = (CICC1851_mainAddrTwo_14 / 2'b10);
  assign CICC1851_mainAddrTwo_14 = ({1'b0,outPixelAddr_value} + CICC1851_mainAddrTwo_15);
  assign CICC1851_mainAddrTwo_16 = {1'b0,1'b1};
  assign CICC1851_mainAddrTwo_15 = {11'd0, CICC1851_mainAddrTwo_16};
  assign CICC1851_counterAddrOne_11 = (CICC1851_counterAddrOne_12 / 2'b10);
  assign CICC1851_counterAddrOne_12 = ({1'b0,outPixelAddr_value} + CICC1851_counterAddrOne_13);
  assign CICC1851_counterAddrOne_14 = {1'b0,1'b1};
  assign CICC1851_counterAddrOne_13 = {11'd0, CICC1851_counterAddrOne_14};
  assign CICC1851_controls_twiceMode_2 = 1'b1;
  assign CICC1851_mainAddrTwo_17 = (CICC1851_mainAddrTwo_18 / 2'b10);
  assign CICC1851_mainAddrTwo_18 = (outPixelAddr_value - 12'h003);
  assign CICC1851_counterAddrOne_15 = (CICC1851_counterAddrOne_16 / 2'b10);
  assign CICC1851_counterAddrOne_16 = (outPixelAddr_value - 12'h003);
  assign CICC1851_mainAddrOne_13 = (CICC1851_mainAddrOne_14 / 2'b10);
  assign CICC1851_mainAddrOne_14 = (outPixelAddr_value - 12'h003);
  assign CICC1851_counterAddrTwo_11 = (CICC1851_counterAddrTwo_12 / 2'b10);
  assign CICC1851_counterAddrTwo_12 = (outPixelAddr_value - 12'h003);
  assign CICC1851_mainAddrOne_15 = (CICC1851_mainAddrOne_16 / 2'b10);
  assign CICC1851_mainAddrOne_16 = ({1'b0,outPixelAddr_value} + CICC1851_mainAddrOne_17);
  assign CICC1851_mainAddrOne_18 = {1'b0,1'b1};
  assign CICC1851_mainAddrOne_17 = {11'd0, CICC1851_mainAddrOne_18};
  assign CICC1851_counterAddrTwo_13 = (CICC1851_counterAddrTwo_14 / 2'b10);
  assign CICC1851_counterAddrTwo_14 = ({1'b0,outPixelAddr_value} + CICC1851_counterAddrTwo_15);
  assign CICC1851_counterAddrTwo_16 = {1'b0,1'b1};
  assign CICC1851_counterAddrTwo_15 = {11'd0, CICC1851_counterAddrTwo_16};
  assign CICC1851_lineBufferOne_port = passPixels_payload_pixel;
  assign CICC1851_lineBufferOne_port_1 = (passPixels_fire_6 && (bufferSwitch == 2'b00));
  assign CICC1851_lineBufferTwo_port = passPixels_payload_pixel;
  assign CICC1851_lineBufferTwo_port_1 = (passPixels_fire_8 && (bufferSwitch == 2'b10));
  assign CICC1851_lineBufferOdd_port = passPixels_payload_pixel;
  assign CICC1851_lineBufferOdd_port_1 = (passPixels_fire_7 && (bufferSwitch == 2'b01));
  always @(posedge clk) begin
    if(CICC1851_lineBufferOne_port_1) begin
      lineBufferOne[bufferWAddr_value] <= CICC1851_lineBufferOne_port;
    end
  end

  always @(posedge clk) begin
    if(mainAddrOneStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferOne_port1 <= lineBufferOne[mainAddrOneStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(counterAddrOneStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferOne_port2 <= lineBufferOne[counterAddrOneStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(CICC1851_lineBufferTwo_port_1) begin
      lineBufferTwo[bufferWAddr_value] <= CICC1851_lineBufferTwo_port;
    end
  end

  always @(posedge clk) begin
    if(mainAddrTwoStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferTwo_port1 <= lineBufferTwo[mainAddrTwoStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(counterAddrTwoStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferTwo_port2 <= lineBufferTwo[counterAddrTwoStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(CICC1851_lineBufferOdd_port_1) begin
      lineBufferOdd[bufferWAddr_value] <= CICC1851_lineBufferOdd_port;
    end
  end

  always @(posedge clk) begin
    if(oddAddrStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferOdd_port1 <= lineBufferOdd[oddAddrStream_s2mPipe_m2sPipe_payload];
    end
  end

  StreamFork_2 diffStage_controlPipe_fork (
    .io_input_valid                      (diffStage_controlPipe_valid                                     ), //i
    .io_input_ready                      (diffStage_controlPipe_fork_io_input_ready                       ), //o
    .io_input_payload_frameStart         (diffStage_controlPipe_payload_frameStart                        ), //i
    .io_input_payload_rowEnd             (diffStage_controlPipe_payload_rowEnd                            ), //i
    .io_input_payload_passMode           (diffStage_controlPipe_payload_passMode                          ), //i
    .io_input_payload_passValid          (diffStage_controlPipe_payload_passValid                         ), //i
    .io_input_payload_onceMode           (diffStage_controlPipe_payload_onceMode[2:0]                     ), //i
    .io_input_payload_onceValid          (diffStage_controlPipe_payload_onceValid                         ), //i
    .io_input_payload_mainCompare        (diffStage_controlPipe_payload_mainCompare                       ), //i
    .io_input_payload_counterCompare     (diffStage_controlPipe_payload_counterCompare                    ), //i
    .io_input_payload_mainDiff           (diffStage_controlPipe_payload_mainDiff[7:0]                     ), //i
    .io_input_payload_counterDiff        (diffStage_controlPipe_payload_counterDiff[7:0]                  ), //i
    .io_input_payload_twiceCompValid     (diffStage_controlPipe_payload_twiceCompValid                    ), //i
    .io_input_payload_twiceMode          (diffStage_controlPipe_payload_twiceMode[2:0]                    ), //i
    .io_input_payload_inpValidFlag       (diffStage_controlPipe_payload_inpValidFlag                      ), //i
    .io_input_payload_oddValid           (diffStage_controlPipe_payload_oddValid                          ), //i
    .io_outputs_0_valid                  (diffStage_controlPipe_fork_io_outputs_0_valid                   ), //o
    .io_outputs_0_ready                  (diffStage_controlPipe_fork_io_outputs_0_translated_ready        ), //i
    .io_outputs_0_payload_frameStart     (diffStage_controlPipe_fork_io_outputs_0_payload_frameStart      ), //o
    .io_outputs_0_payload_rowEnd         (diffStage_controlPipe_fork_io_outputs_0_payload_rowEnd          ), //o
    .io_outputs_0_payload_passMode       (diffStage_controlPipe_fork_io_outputs_0_payload_passMode        ), //o
    .io_outputs_0_payload_passValid      (diffStage_controlPipe_fork_io_outputs_0_payload_passValid       ), //o
    .io_outputs_0_payload_onceMode       (diffStage_controlPipe_fork_io_outputs_0_payload_onceMode[2:0]   ), //o
    .io_outputs_0_payload_onceValid      (diffStage_controlPipe_fork_io_outputs_0_payload_onceValid       ), //o
    .io_outputs_0_payload_mainCompare    (diffStage_controlPipe_fork_io_outputs_0_payload_mainCompare     ), //o
    .io_outputs_0_payload_counterCompare (diffStage_controlPipe_fork_io_outputs_0_payload_counterCompare  ), //o
    .io_outputs_0_payload_mainDiff       (diffStage_controlPipe_fork_io_outputs_0_payload_mainDiff[7:0]   ), //o
    .io_outputs_0_payload_counterDiff    (diffStage_controlPipe_fork_io_outputs_0_payload_counterDiff[7:0]), //o
    .io_outputs_0_payload_twiceCompValid (diffStage_controlPipe_fork_io_outputs_0_payload_twiceCompValid  ), //o
    .io_outputs_0_payload_twiceMode      (diffStage_controlPipe_fork_io_outputs_0_payload_twiceMode[2:0]  ), //o
    .io_outputs_0_payload_inpValidFlag   (diffStage_controlPipe_fork_io_outputs_0_payload_inpValidFlag    ), //o
    .io_outputs_0_payload_oddValid       (diffStage_controlPipe_fork_io_outputs_0_payload_oddValid        ), //o
    .io_outputs_1_valid                  (diffStage_controlPipe_fork_io_outputs_1_valid                   ), //o
    .io_outputs_1_ready                  (resultStage_pixelStream_ready                                   ), //i
    .io_outputs_1_payload_frameStart     (diffStage_controlPipe_fork_io_outputs_1_payload_frameStart      ), //o
    .io_outputs_1_payload_rowEnd         (diffStage_controlPipe_fork_io_outputs_1_payload_rowEnd          ), //o
    .io_outputs_1_payload_passMode       (diffStage_controlPipe_fork_io_outputs_1_payload_passMode        ), //o
    .io_outputs_1_payload_passValid      (diffStage_controlPipe_fork_io_outputs_1_payload_passValid       ), //o
    .io_outputs_1_payload_onceMode       (diffStage_controlPipe_fork_io_outputs_1_payload_onceMode[2:0]   ), //o
    .io_outputs_1_payload_onceValid      (diffStage_controlPipe_fork_io_outputs_1_payload_onceValid       ), //o
    .io_outputs_1_payload_mainCompare    (diffStage_controlPipe_fork_io_outputs_1_payload_mainCompare     ), //o
    .io_outputs_1_payload_counterCompare (diffStage_controlPipe_fork_io_outputs_1_payload_counterCompare  ), //o
    .io_outputs_1_payload_mainDiff       (diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff[7:0]   ), //o
    .io_outputs_1_payload_counterDiff    (diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff[7:0]), //o
    .io_outputs_1_payload_twiceCompValid (diffStage_controlPipe_fork_io_outputs_1_payload_twiceCompValid  ), //o
    .io_outputs_1_payload_twiceMode      (diffStage_controlPipe_fork_io_outputs_1_payload_twiceMode[2:0]  ), //o
    .io_outputs_1_payload_inpValidFlag   (diffStage_controlPipe_fork_io_outputs_1_payload_inpValidFlag    ), //o
    .io_outputs_1_payload_oddValid       (diffStage_controlPipe_fork_io_outputs_1_payload_oddValid        )  //o
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_1_BOOT : controlStateMachine_stateReg_string = "BOOT ";
      controlStateMachine_enumDef_1_HOLD : controlStateMachine_stateReg_string = "HOLD ";
      controlStateMachine_enumDef_1_PASS : controlStateMachine_stateReg_string = "PASS ";
      controlStateMachine_enumDef_1_ONCE : controlStateMachine_stateReg_string = "ONCE ";
      controlStateMachine_enumDef_1_TWICE : controlStateMachine_stateReg_string = "TWICE";
      default : controlStateMachine_stateReg_string = "?????";
    endcase
  end
  always @(*) begin
    case(controlStateMachine_stateNext)
      controlStateMachine_enumDef_1_BOOT : controlStateMachine_stateNext_string = "BOOT ";
      controlStateMachine_enumDef_1_HOLD : controlStateMachine_stateNext_string = "HOLD ";
      controlStateMachine_enumDef_1_PASS : controlStateMachine_stateNext_string = "PASS ";
      controlStateMachine_enumDef_1_ONCE : controlStateMachine_stateNext_string = "ONCE ";
      controlStateMachine_enumDef_1_TWICE : controlStateMachine_stateNext_string = "TWICE";
      default : controlStateMachine_stateNext_string = "?????";
    endcase
  end
  `endif

  always @(*) begin
    pixelsIn_ready = 1'b0;
    pixelsIn_ready = (! pixelsIn_rValid);
  end

  always @(*) begin
    pixelsOut_valid = 1'b0;
    pixelsOut_valid = pixelsStream_s2mPipe_m2sPipe_valid;
  end

  always @(*) begin
    pixelsOut_payload_pixel = 8'h0;
    pixelsOut_payload_pixel = pixelsStream_s2mPipe_m2sPipe_payload_pixel;
  end

  always @(*) begin
    pixelsOut_payload_frameStart = 1'b0;
    pixelsOut_payload_frameStart = pixelsStream_s2mPipe_m2sPipe_payload_frameStart;
  end

  always @(*) begin
    pixelsOut_payload_rowEnd = 1'b0;
    pixelsOut_payload_rowEnd = pixelsStream_s2mPipe_m2sPipe_payload_rowEnd;
  end

  always @(*) begin
    pixelsOut_payload_inpValid = 1'b0;
    pixelsOut_payload_inpValid = pixelsStream_s2mPipe_m2sPipe_payload_inpValid;
  end

  always @(*) begin
    startOut = 1'b0;
    startOut = slaveStart;
  end

  always @(*) begin
    inpTwoDoneOut = 1'b0;
    inpTwoDoneOut = inpTwoDone;
  end

  assign when_SuperResolutionPart2_l40 = (inpThreeDoneIn || (startIn && (! startIn_regNext)));
  assign when_SuperResolutionPart2_l43 = (! startIn);
  assign when_SuperResolutionPart2_l46 = (startIn && (! readDone));
  assign when_SuperResolutionPart2_l46_1 = (! startIn);
  assign pixelsIn_fire = (pixelsIn_valid && pixelsIn_ready);
  assign when_SuperResolutionPart2_l49 = ((! inpThreeDoneIn) && pixelsIn_fire);
  assign when_SuperResolutionPart2_l49_1 = (inpThreeDoneIn || (! startIn));
  assign when_SuperResolutionPart2_l64 = (! startIn);
  assign when_SuperResolutionPart2_l67 = (! startIn);
  always @(*) begin
    bufferRowCount_willIncrement = 1'b0;
    if(when_SuperResolutionPart2_l185) begin
      if(!bufferReachFinalRow) begin
        bufferRowCount_willIncrement = 1'b1;
      end
    end
  end

  always @(*) begin
    bufferRowCount_willClear = 1'b0;
    if(when_SuperResolutionPart2_l185) begin
      if(bufferReachFinalRow) begin
        bufferRowCount_willClear = 1'b1;
      end
    end
  end

  assign bufferRowCount_willOverflowIfInc = (bufferRowCount_value == 11'h438);
  assign bufferRowCount_willOverflow = (bufferRowCount_willOverflowIfInc && bufferRowCount_willIncrement);
  always @(*) begin
    if(bufferRowCount_willOverflow) begin
      bufferRowCount_valueNext = 11'h0;
    end else begin
      bufferRowCount_valueNext = (bufferRowCount_value + CICC1851_bufferRowCount_valueNext);
    end
    if(bufferRowCount_willClear) begin
      bufferRowCount_valueNext = 11'h0;
    end
  end

  assign when_SuperResolutionPart2_l76 = ((startIn && (! holdBuffer)) && (! writeDone));
  assign when_SuperResolutionPart2_l76_1 = (((! startIn) || holdBuffer) || writeDone);
  assign when_SuperResolutionPart2_l82 = (! startRead);
  always @(*) begin
    bufferWAddr_willIncrement = 1'b0;
    if(passPixels_fire_9) begin
      if(!passPixels_payload_rowEnd) begin
        bufferWAddr_willIncrement = 1'b1;
      end
    end
  end

  always @(*) begin
    bufferWAddr_willClear = 1'b0;
    if(passPixels_fire_9) begin
      if(passPixels_payload_rowEnd) begin
        bufferWAddr_willClear = 1'b1;
      end
    end
  end

  assign bufferWAddr_willOverflowIfInc = (bufferWAddr_value == 11'h77f);
  assign bufferWAddr_willOverflow = (bufferWAddr_willOverflowIfInc && bufferWAddr_willIncrement);
  always @(*) begin
    if(bufferWAddr_willOverflow) begin
      bufferWAddr_valueNext = 11'h0;
    end else begin
      bufferWAddr_valueNext = (bufferWAddr_value + CICC1851_bufferWAddr_valueNext);
    end
    if(bufferWAddr_willClear) begin
      bufferWAddr_valueNext = 11'h0;
    end
  end

  always @(*) begin
    outPixelAddr_willIncrement = 1'b0;
    if(when_SuperResolutionPart2_l761) begin
      if(controlStream_fire_7) begin
        if(!outReachRowEnd) begin
          outPixelAddr_willIncrement = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    outPixelAddr_willClear = 1'b0;
    if(when_SuperResolutionPart2_l761) begin
      if(controlStream_fire_7) begin
        if(outReachRowEnd) begin
          outPixelAddr_willClear = 1'b1;
        end
      end
    end
  end

  assign outPixelAddr_willOverflowIfInc = (outPixelAddr_value == 12'heff);
  assign outPixelAddr_willOverflow = (outPixelAddr_willOverflowIfInc && outPixelAddr_willIncrement);
  always @(*) begin
    if(outPixelAddr_willOverflow) begin
      outPixelAddr_valueNext = 12'h0;
    end else begin
      outPixelAddr_valueNext = (outPixelAddr_value + CICC1851_outPixelAddr_valueNext);
    end
    if(outPixelAddr_willClear) begin
      outPixelAddr_valueNext = 12'h0;
    end
  end

  always @(*) begin
    outRowCount_willIncrement = 1'b0;
    if(when_SuperResolutionPart2_l761) begin
      if(when_SuperResolutionPart2_l766) begin
        if(!outReachFinalRow) begin
          outRowCount_willIncrement = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    outRowCount_willClear = 1'b0;
    if(when_SuperResolutionPart2_l761) begin
      if(when_SuperResolutionPart2_l766) begin
        if(outReachFinalRow) begin
          outRowCount_willClear = 1'b1;
        end
      end
    end
  end

  assign outRowCount_willOverflowIfInc = (outRowCount_value == 12'h870);
  assign outRowCount_willOverflow = (outRowCount_willOverflowIfInc && outRowCount_willIncrement);
  always @(*) begin
    if(outRowCount_willOverflow) begin
      outRowCount_valueNext = 12'h0;
    end else begin
      outRowCount_valueNext = (outRowCount_value + CICC1851_outRowCount_valueNext);
    end
    if(outRowCount_willClear) begin
      outRowCount_valueNext = 12'h0;
    end
  end

  always @(*) begin
    alreadySendRow_willIncrement = 1'b0;
    if(pixelsOut_fire_2) begin
      if(alreadyReachRowEnd) begin
        if(!alreadyReachFinalRow) begin
          alreadySendRow_willIncrement = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    alreadySendRow_willClear = 1'b0;
    if(pixelsOut_fire_2) begin
      if(alreadyReachRowEnd) begin
        if(alreadyReachFinalRow) begin
          alreadySendRow_willClear = 1'b1;
        end
      end
    end
  end

  assign alreadySendRow_willOverflowIfInc = (alreadySendRow_value == 12'h870);
  assign alreadySendRow_willOverflow = (alreadySendRow_willOverflowIfInc && alreadySendRow_willIncrement);
  always @(*) begin
    if(alreadySendRow_willOverflow) begin
      alreadySendRow_valueNext = 12'h0;
    end else begin
      alreadySendRow_valueNext = (alreadySendRow_value + CICC1851_alreadySendRow_valueNext);
    end
    if(alreadySendRow_willClear) begin
      alreadySendRow_valueNext = 12'h0;
    end
  end

  always @(*) begin
    alreadySendCountInRow_willIncrement = 1'b0;
    if(pixelsOut_fire_2) begin
      if(!alreadyReachRowEnd) begin
        alreadySendCountInRow_willIncrement = 1'b1;
      end
    end
  end

  always @(*) begin
    alreadySendCountInRow_willClear = 1'b0;
    if(pixelsOut_fire_2) begin
      if(alreadyReachRowEnd) begin
        alreadySendCountInRow_willClear = 1'b1;
      end
    end
  end

  assign alreadySendCountInRow_willOverflowIfInc = (alreadySendCountInRow_value == 12'heff);
  assign alreadySendCountInRow_willOverflow = (alreadySendCountInRow_willOverflowIfInc && alreadySendCountInRow_willIncrement);
  always @(*) begin
    if(alreadySendCountInRow_willOverflow) begin
      alreadySendCountInRow_valueNext = 12'h0;
    end else begin
      alreadySendCountInRow_valueNext = (alreadySendCountInRow_value + CICC1851_alreadySendCountInRow_valueNext);
    end
    if(alreadySendCountInRow_willClear) begin
      alreadySendCountInRow_valueNext = 12'h0;
    end
  end

  assign when_SuperResolutionPart2_l106 = (((! startIn) && startIn_regNext_1) || inpTwoDone);
  assign when_SuperResolutionPart2_l108 = (((! startIn) && startIn_regNext_2) || inpTwoDone);
  assign when_SuperResolutionPart2_l109 = (((! startIn) && startIn_regNext_3) || inpTwoDone);
  assign when_SuperResolutionPart2_l110 = (((! startIn) && startIn_regNext_4) || inpTwoDone);
  assign when_SuperResolutionPart2_l111 = (((! startIn) && startIn_regNext_5) || inpTwoDone);
  assign when_SuperResolutionPart2_l113 = (((! startIn) && startIn_regNext_6) || inpTwoDone);
  assign when_SuperResolutionPart2_l114 = (((! startIn) && startIn_regNext_7) || inpTwoDone);
  assign when_SuperResolutionPart2_l115 = (((! startIn) && startIn_regNext_8) || inpTwoDone);
  assign when_SuperResolutionPart2_l116 = (((! startIn) && startIn_regNext_9) || inpTwoDone);
  assign when_SuperResolutionPart2_l120 = (((! startIn) && startIn_regNext_10) || inpTwoDone);
  assign when_SuperResolutionPart2_l121 = (((! startIn) && startIn_regNext_11) || inpTwoDone);
  assign when_SuperResolutionPart2_l122 = (((! startIn) && startIn_regNext_12) || inpTwoDone);
  assign when_SuperResolutionPart2_l123 = (((! startIn) && startIn_regNext_13) || inpTwoDone);
  assign when_SuperResolutionPart2_l124 = (((! startIn) && startIn_regNext_14) || inpTwoDone);
  assign when_SuperResolutionPart2_l125 = (((! startIn) && startIn_regNext_15) || inpTwoDone);
  assign when_SuperResolutionPart2_l126 = (((! startIn) && startIn_regNext_16) || inpTwoDone);
  assign when_SuperResolutionPart2_l134 = (! startRead);
  always @(*) begin
    mainAddrOne = CICC1851_mainAddrOne[10:0];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_1_HOLD : begin
      end
      controlStateMachine_enumDef_1_PASS : begin
        if(!twoInFourOutRow) begin
          if(oneInFourOutRow) begin
            if(nextRowBuffer) begin
              if(twoInFourOutPixelAddr) begin
                mainAddrOne = CICC1851_mainAddrOne_1[10:0];
              end
            end
          end
        end
      end
      controlStateMachine_enumDef_1_ONCE : begin
        if(threeInFourOutRow) begin
          if(twoInFourOutPixelAddr) begin
            mainAddrOne = CICC1851_mainAddrOne_3[10:0];
          end
        end else begin
          if(nextRowBuffer) begin
            mainAddrOne = CICC1851_mainAddrOne_5[10:0];
          end
        end
      end
      controlStateMachine_enumDef_1_TWICE : begin
        if(outReachFinalRow) begin
          if(nextRowBuffer) begin
            if(outReachRowEnd) begin
              mainAddrOne = CICC1851_mainAddrOne_7[10:0];
            end else begin
              mainAddrOne = CICC1851_mainAddrOne_9[10:0];
            end
          end
        end else begin
          if(nextRowBuffer) begin
            mainAddrOne = CICC1851_mainAddrOne_11[10:0];
          end else begin
            if(outReachRowEnd) begin
              mainAddrOne = CICC1851_mainAddrOne_13[10:0];
            end else begin
              mainAddrOne = CICC1851_mainAddrOne_15[10:0];
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    counterAddrOne = CICC1851_counterAddrOne[10:0];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_1_HOLD : begin
      end
      controlStateMachine_enumDef_1_PASS : begin
      end
      controlStateMachine_enumDef_1_ONCE : begin
        if(!threeInFourOutRow) begin
          if(nextRowBuffer) begin
            if(outReachRowEnd) begin
              counterAddrOne = CICC1851_counterAddrOne_1[10:0];
            end else begin
              counterAddrOne = CICC1851_counterAddrOne_3[10:0];
            end
          end
        end
      end
      controlStateMachine_enumDef_1_TWICE : begin
        if(outReachFinalRow) begin
          if(nextRowBuffer) begin
            if(!outReachRowEnd) begin
              counterAddrOne = CICC1851_counterAddrOne_5[10:0];
            end
          end
        end else begin
          if(nextRowBuffer) begin
            if(outReachRowEnd) begin
              counterAddrOne = CICC1851_counterAddrOne_9[10:0];
            end else begin
              counterAddrOne = CICC1851_counterAddrOne_11[10:0];
            end
          end else begin
            counterAddrOne = CICC1851_counterAddrOne_15[10:0];
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    mainAddrTwo = CICC1851_mainAddrTwo[10:0];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_1_HOLD : begin
      end
      controlStateMachine_enumDef_1_PASS : begin
        if(!twoInFourOutRow) begin
          if(oneInFourOutRow) begin
            if(!nextRowBuffer) begin
              if(twoInFourOutPixelAddr) begin
                mainAddrTwo = CICC1851_mainAddrTwo_1[10:0];
              end
            end
          end
        end
      end
      controlStateMachine_enumDef_1_ONCE : begin
        if(threeInFourOutRow) begin
          if(twoInFourOutPixelAddr) begin
            mainAddrTwo = CICC1851_mainAddrTwo_3[10:0];
          end
        end else begin
          if(!nextRowBuffer) begin
            mainAddrTwo = CICC1851_mainAddrTwo_5[10:0];
          end
        end
      end
      controlStateMachine_enumDef_1_TWICE : begin
        if(outReachFinalRow) begin
          if(!nextRowBuffer) begin
            if(outReachRowEnd) begin
              mainAddrTwo = CICC1851_mainAddrTwo_7[10:0];
            end else begin
              mainAddrTwo = CICC1851_mainAddrTwo_9[10:0];
            end
          end
        end else begin
          if(nextRowBuffer) begin
            if(outReachRowEnd) begin
              mainAddrTwo = CICC1851_mainAddrTwo_11[10:0];
            end else begin
              mainAddrTwo = CICC1851_mainAddrTwo_13[10:0];
            end
          end else begin
            mainAddrTwo = CICC1851_mainAddrTwo_17[10:0];
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    counterAddrTwo = CICC1851_counterAddrTwo[10:0];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_1_HOLD : begin
      end
      controlStateMachine_enumDef_1_PASS : begin
      end
      controlStateMachine_enumDef_1_ONCE : begin
        if(!threeInFourOutRow) begin
          if(!nextRowBuffer) begin
            if(outReachRowEnd) begin
              counterAddrTwo = CICC1851_counterAddrTwo_1[10:0];
            end else begin
              counterAddrTwo = CICC1851_counterAddrTwo_3[10:0];
            end
          end
        end
      end
      controlStateMachine_enumDef_1_TWICE : begin
        if(outReachFinalRow) begin
          if(!nextRowBuffer) begin
            if(!outReachRowEnd) begin
              counterAddrTwo = CICC1851_counterAddrTwo_5[10:0];
            end
          end
        end else begin
          if(nextRowBuffer) begin
            counterAddrTwo = CICC1851_counterAddrTwo_9[10:0];
          end else begin
            if(outReachRowEnd) begin
              counterAddrTwo = CICC1851_counterAddrTwo_11[10:0];
            end else begin
              counterAddrTwo = CICC1851_counterAddrTwo_13[10:0];
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign oddAddr = CICC1851_oddAddr[10:0];
  assign validStream_valid = 1'b1;
  assign CICC1851_controls_frameStart = 32'h0;
  always @(*) begin
    controls_frameStart = CICC1851_controls_frameStart[0];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_1_HOLD : begin
      end
      controlStateMachine_enumDef_1_PASS : begin
        if(frameStart) begin
          controls_frameStart = 1'b1;
        end
      end
      controlStateMachine_enumDef_1_ONCE : begin
      end
      controlStateMachine_enumDef_1_TWICE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_rowEnd = CICC1851_controls_frameStart[1];
    if(when_SuperResolutionPart2_l761) begin
      if(outReachRowEnd) begin
        controls_rowEnd = 1'b1;
      end
    end
  end

  always @(*) begin
    controls_passMode = CICC1851_controls_frameStart[2];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_1_HOLD : begin
      end
      controlStateMachine_enumDef_1_PASS : begin
        if(twoInFourOutRow) begin
          if(!when_SuperResolutionPart2_l609) begin
            if(nextRowBuffer) begin
              controls_passMode = 1'b0;
            end else begin
              controls_passMode = 1'b1;
            end
          end
        end else begin
          if(oneInFourOutRow) begin
            if(nextRowBuffer) begin
              controls_passMode = 1'b0;
            end else begin
              controls_passMode = 1'b1;
            end
          end else begin
            if(nextRowBuffer) begin
              controls_passMode = 1'b0;
            end else begin
              controls_passMode = 1'b1;
            end
          end
        end
      end
      controlStateMachine_enumDef_1_ONCE : begin
      end
      controlStateMachine_enumDef_1_TWICE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_passValid = CICC1851_controls_frameStart[3];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_1_HOLD : begin
      end
      controlStateMachine_enumDef_1_PASS : begin
        if(twoInFourOutRow) begin
          if(!when_SuperResolutionPart2_l609) begin
            controls_passValid = 1'b1;
          end
        end else begin
          if(oneInFourOutRow) begin
            controls_passValid = 1'b1;
          end else begin
            controls_passValid = 1'b1;
          end
        end
      end
      controlStateMachine_enumDef_1_ONCE : begin
      end
      controlStateMachine_enumDef_1_TWICE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_onceMode = CICC1851_controls_frameStart[6 : 4];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_1_HOLD : begin
      end
      controlStateMachine_enumDef_1_PASS : begin
      end
      controlStateMachine_enumDef_1_ONCE : begin
        if(threeInFourOutRow) begin
          if(outReachFinalRow) begin
            if(nextRowBuffer) begin
              controls_onceMode = 3'b100;
            end else begin
              controls_onceMode = 3'b101;
            end
          end else begin
            if(nextRowBuffer) begin
              controls_onceMode = {1'd0, CICC1851_controls_onceMode};
            end else begin
              controls_onceMode = {1'd0, CICC1851_controls_onceMode_1};
            end
          end
        end else begin
          if(nextRowBuffer) begin
            controls_onceMode = 3'b000;
          end else begin
            controls_onceMode = {2'd0, CICC1851_controls_onceMode_2};
          end
        end
      end
      controlStateMachine_enumDef_1_TWICE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_onceValid = CICC1851_controls_frameStart[7];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_1_HOLD : begin
      end
      controlStateMachine_enumDef_1_PASS : begin
      end
      controlStateMachine_enumDef_1_ONCE : begin
        controls_onceValid = 1'b1;
      end
      controlStateMachine_enumDef_1_TWICE : begin
      end
      default : begin
      end
    endcase
  end

  assign controls_mainCompare = CICC1851_controls_frameStart[8];
  assign controls_counterCompare = CICC1851_controls_frameStart[9];
  assign controls_mainDiff = CICC1851_controls_frameStart[17 : 10];
  assign controls_counterDiff = CICC1851_controls_frameStart[25 : 18];
  always @(*) begin
    controls_twiceCompValid = CICC1851_controls_frameStart[26];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_1_HOLD : begin
      end
      controlStateMachine_enumDef_1_PASS : begin
      end
      controlStateMachine_enumDef_1_ONCE : begin
      end
      controlStateMachine_enumDef_1_TWICE : begin
        controls_twiceCompValid = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_twiceMode = CICC1851_controls_frameStart[29 : 27];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_1_HOLD : begin
      end
      controlStateMachine_enumDef_1_PASS : begin
      end
      controlStateMachine_enumDef_1_ONCE : begin
      end
      controlStateMachine_enumDef_1_TWICE : begin
        if(outReachFinalRow) begin
          if(nextRowBuffer) begin
            if(outReachRowEnd) begin
              controls_twiceMode = 3'b100;
            end else begin
              controls_twiceMode = 3'b101;
            end
          end else begin
            if(outReachRowEnd) begin
              controls_twiceMode = {1'd0, CICC1851_controls_twiceMode};
            end else begin
              controls_twiceMode = {1'd0, CICC1851_controls_twiceMode_1};
            end
          end
        end else begin
          if(nextRowBuffer) begin
            controls_twiceMode = 3'b000;
          end else begin
            controls_twiceMode = {2'd0, CICC1851_controls_twiceMode_2};
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_inpValidFlag = CICC1851_controls_frameStart[30];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_1_HOLD : begin
        controls_inpValidFlag = 1'b1;
      end
      controlStateMachine_enumDef_1_PASS : begin
        controls_inpValidFlag = 1'b1;
      end
      controlStateMachine_enumDef_1_ONCE : begin
        controls_inpValidFlag = 1'b1;
      end
      controlStateMachine_enumDef_1_TWICE : begin
        controls_inpValidFlag = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_oddValid = CICC1851_controls_frameStart[31];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_1_HOLD : begin
      end
      controlStateMachine_enumDef_1_PASS : begin
        if(twoInFourOutRow) begin
          if(when_SuperResolutionPart2_l609) begin
            controls_oddValid = 1'b1;
          end
        end
      end
      controlStateMachine_enumDef_1_ONCE : begin
      end
      controlStateMachine_enumDef_1_TWICE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    validStream_ready = (controlStream_ready && startRead);
    validStream_ready = (mainAddrOneStream_ready && startRead);
    validStream_ready = (counterAddrOneStream_ready && startRead);
    validStream_ready = (mainAddrTwoStream_ready && startRead);
    validStream_ready = (counterAddrTwoStream_ready && startRead);
    validStream_ready = (oddAddrStream_ready && startRead);
  end

  assign controlStream_valid = (validStream_valid && startRead);
  assign controlStream_payload_frameStart = controls_frameStart;
  assign controlStream_payload_rowEnd = controls_rowEnd;
  assign controlStream_payload_passMode = controls_passMode;
  assign controlStream_payload_passValid = controls_passValid;
  assign controlStream_payload_onceMode = controls_onceMode;
  assign controlStream_payload_onceValid = controls_onceValid;
  assign controlStream_payload_mainCompare = controls_mainCompare;
  assign controlStream_payload_counterCompare = controls_counterCompare;
  assign controlStream_payload_mainDiff = controls_mainDiff;
  assign controlStream_payload_counterDiff = controls_counterDiff;
  assign controlStream_payload_twiceCompValid = controls_twiceCompValid;
  assign controlStream_payload_twiceMode = controls_twiceMode;
  assign controlStream_payload_inpValidFlag = controls_inpValidFlag;
  assign controlStream_payload_oddValid = controls_oddValid;
  assign mainAddrOneStream_valid = (validStream_valid && startRead);
  assign mainAddrOneStream_payload = mainAddrOne;
  assign counterAddrOneStream_valid = (validStream_valid && startRead);
  assign counterAddrOneStream_payload = counterAddrOne;
  assign mainAddrTwoStream_valid = (validStream_valid && startRead);
  assign mainAddrTwoStream_payload = mainAddrTwo;
  assign counterAddrTwoStream_valid = (validStream_valid && startRead);
  assign counterAddrTwoStream_payload = counterAddrTwo;
  assign oddAddrStream_valid = (validStream_valid && startRead);
  assign oddAddrStream_payload = oddAddr;
  assign pixelsIn_s2mPipe_valid = (pixelsIn_valid || pixelsIn_rValid);
  assign pixelsIn_s2mPipe_payload_pixel = (pixelsIn_rValid ? pixelsIn_rData_pixel : pixelsIn_payload_pixel);
  assign pixelsIn_s2mPipe_payload_frameStart = (pixelsIn_rValid ? pixelsIn_rData_frameStart : pixelsIn_payload_frameStart);
  assign pixelsIn_s2mPipe_payload_rowEnd = (pixelsIn_rValid ? pixelsIn_rData_rowEnd : pixelsIn_payload_rowEnd);
  always @(*) begin
    pixelsIn_s2mPipe_ready = pixelsIn_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368) begin
      pixelsIn_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368 = (! pixelsIn_s2mPipe_m2sPipe_valid);
  assign pixelsIn_s2mPipe_m2sPipe_valid = pixelsIn_s2mPipe_rValid;
  assign pixelsIn_s2mPipe_m2sPipe_payload_pixel = pixelsIn_s2mPipe_rData_pixel;
  assign pixelsIn_s2mPipe_m2sPipe_payload_frameStart = pixelsIn_s2mPipe_rData_frameStart;
  assign pixelsIn_s2mPipe_m2sPipe_payload_rowEnd = pixelsIn_s2mPipe_rData_rowEnd;
  assign passPixels_valid = (pixelsIn_s2mPipe_m2sPipe_valid && bufferEnable);
  assign pixelsIn_s2mPipe_m2sPipe_ready = (passPixels_ready && bufferEnable);
  assign passPixels_payload_pixel = pixelsIn_s2mPipe_m2sPipe_payload_pixel;
  assign passPixels_payload_frameStart = pixelsIn_s2mPipe_m2sPipe_payload_frameStart;
  assign passPixels_payload_rowEnd = pixelsIn_s2mPipe_m2sPipe_payload_rowEnd;
  assign passPixels_ready = 1'b1;
  assign passPixels_fire = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart2_l181 = ((CICC1851_when_SuperResolutionPart2_l181 == CICC1851_when_SuperResolutionPart2_l181_1) && passPixels_fire);
  assign passPixels_fire_1 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart2_l182 = (((CICC1851_when_SuperResolutionPart2_l182 == CICC1851_when_SuperResolutionPart2_l182_1) && bufferReachRowEnd) && passPixels_fire_1);
  assign passPixels_fire_2 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart2_l185 = (passPixels_payload_rowEnd && passPixels_fire_2);
  assign when_SuperResolutionPart2_l195 = (CICC1851_when_SuperResolutionPart2_l195 == 11'h0);
  assign passPixels_fire_3 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart2_l200 = (passPixels_payload_rowEnd && passPixels_fire_3);
  assign when_SuperResolutionPart2_l201 = ((bufferSwitch == 2'b10) || (bufferSwitch == 2'b00));
  assign passPixels_fire_4 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart2_l207 = (((bufferRowCount_value != 11'h0) && passPixels_payload_rowEnd) && passPixels_fire_4);
  assign when_SuperResolutionPart2_l208 = (bufferSwitch != 2'b01);
  assign when_SuperResolutionPart2_l212 = (bufferReachFinalRow && bufferReachRowEnd);
  assign controlStream_fire = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart2_l218 = (((CICC1851_when_SuperResolutionPart2_l218 == 12'h003) && controlStream_payload_rowEnd) && controlStream_fire);
  assign when_SuperResolutionPart2_l220 = 1'b1;
  assign passPixels_fire_5 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart2_l224 = (passPixels_payload_frameStart && passPixels_fire_5);
  assign pixelsOut_fire = (pixelsOut_valid && pixelsOut_ready);
  assign when_SuperResolutionPart2_l234 = ((CICC1851_when_SuperResolutionPart2_l234 == CICC1851_when_SuperResolutionPart2_l234_1) && pixelsOut_fire);
  assign pixelsOut_fire_1 = (pixelsOut_valid && pixelsOut_ready);
  assign when_SuperResolutionPart2_l235 = (((CICC1851_when_SuperResolutionPart2_l235 == CICC1851_when_SuperResolutionPart2_l235_1) && alreadyReachRowEnd) && pixelsOut_fire_1);
  assign pixelsOut_fire_2 = (pixelsOut_valid && pixelsOut_ready);
  assign pixelsOut_fire_3 = (pixelsOut_valid && pixelsOut_ready);
  assign when_SuperResolutionPart2_l246 = ((alreadyReachFinalRow && alreadyReachRowEnd) && pixelsOut_fire_3);
  assign passPixels_fire_6 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_7 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_8 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_9 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_10 = (passPixels_valid && passPixels_ready);
  assign controlStream_fire_1 = (controlStream_valid && controlStream_ready);
  assign pushing = (passPixels_fire_10 && (! controlStream_fire_1));
  assign passPixels_fire_11 = (passPixels_valid && passPixels_ready);
  assign controlStream_fire_2 = (controlStream_valid && controlStream_ready);
  assign poping = ((! passPixels_fire_11) && controlStream_fire_2);
  assign passPixels_fire_12 = (passPixels_valid && passPixels_ready);
  assign controlStream_fire_3 = (controlStream_valid && controlStream_ready);
  assign pushAndPoping = (passPixels_fire_12 && controlStream_fire_3);
  assign mainAddrOneStream_ready = (! mainAddrOneStream_rValid);
  assign mainAddrOneStream_s2mPipe_valid = (mainAddrOneStream_valid || mainAddrOneStream_rValid);
  assign mainAddrOneStream_s2mPipe_payload = (mainAddrOneStream_rValid ? mainAddrOneStream_rData : mainAddrOneStream_payload);
  always @(*) begin
    mainAddrOneStream_s2mPipe_ready = mainAddrOneStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_1) begin
      mainAddrOneStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_1 = (! mainAddrOneStream_s2mPipe_m2sPipe_valid);
  assign mainAddrOneStream_s2mPipe_m2sPipe_valid = mainAddrOneStream_s2mPipe_rValid;
  assign mainAddrOneStream_s2mPipe_m2sPipe_payload = mainAddrOneStream_s2mPipe_rData;
  assign mainAddrOneStream_s2mPipe_m2sPipe_ready = ((! CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready) || CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready = CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_mainOnePixelStream_payload = CICC1851_lineBufferOne_port1;
  assign CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_1 = readStage_mainOnePixelStream_ready;
    if(when_Stream_l368_2) begin
      CICC1851_1 = 1'b1;
    end
  end

  assign when_Stream_l368_2 = (! readStage_mainOnePixelStream_valid);
  assign readStage_mainOnePixelStream_valid = CICC1851_readStage_mainOnePixelStream_valid;
  assign readStage_mainOnePixelStream_payload = CICC1851_readStage_mainOnePixelStream_payload_2;
  assign counterAddrOneStream_ready = (! counterAddrOneStream_rValid);
  assign counterAddrOneStream_s2mPipe_valid = (counterAddrOneStream_valid || counterAddrOneStream_rValid);
  assign counterAddrOneStream_s2mPipe_payload = (counterAddrOneStream_rValid ? counterAddrOneStream_rData : counterAddrOneStream_payload);
  always @(*) begin
    counterAddrOneStream_s2mPipe_ready = counterAddrOneStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_3) begin
      counterAddrOneStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_3 = (! counterAddrOneStream_s2mPipe_m2sPipe_valid);
  assign counterAddrOneStream_s2mPipe_m2sPipe_valid = counterAddrOneStream_s2mPipe_rValid;
  assign counterAddrOneStream_s2mPipe_m2sPipe_payload = counterAddrOneStream_s2mPipe_rData;
  assign counterAddrOneStream_s2mPipe_m2sPipe_ready = ((! CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready) || CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready = CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_counterOnePixelStream_payload = CICC1851_lineBufferOne_port2;
  assign CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_2 = readStage_counterOnePixelStream_ready;
    if(when_Stream_l368_4) begin
      CICC1851_2 = 1'b1;
    end
  end

  assign when_Stream_l368_4 = (! readStage_counterOnePixelStream_valid);
  assign readStage_counterOnePixelStream_valid = CICC1851_readStage_counterOnePixelStream_valid;
  assign readStage_counterOnePixelStream_payload = CICC1851_readStage_counterOnePixelStream_payload_2;
  assign mainAddrTwoStream_ready = (! mainAddrTwoStream_rValid);
  assign mainAddrTwoStream_s2mPipe_valid = (mainAddrTwoStream_valid || mainAddrTwoStream_rValid);
  assign mainAddrTwoStream_s2mPipe_payload = (mainAddrTwoStream_rValid ? mainAddrTwoStream_rData : mainAddrTwoStream_payload);
  always @(*) begin
    mainAddrTwoStream_s2mPipe_ready = mainAddrTwoStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_5) begin
      mainAddrTwoStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_5 = (! mainAddrTwoStream_s2mPipe_m2sPipe_valid);
  assign mainAddrTwoStream_s2mPipe_m2sPipe_valid = mainAddrTwoStream_s2mPipe_rValid;
  assign mainAddrTwoStream_s2mPipe_m2sPipe_payload = mainAddrTwoStream_s2mPipe_rData;
  assign mainAddrTwoStream_s2mPipe_m2sPipe_ready = ((! CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready) || CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready = CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_mainTwoPixelStream_payload = CICC1851_lineBufferTwo_port1;
  assign CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_3 = readStage_mainTwoPixelStream_ready;
    if(when_Stream_l368_6) begin
      CICC1851_3 = 1'b1;
    end
  end

  assign when_Stream_l368_6 = (! readStage_mainTwoPixelStream_valid);
  assign readStage_mainTwoPixelStream_valid = CICC1851_readStage_mainTwoPixelStream_valid;
  assign readStage_mainTwoPixelStream_payload = CICC1851_readStage_mainTwoPixelStream_payload_2;
  assign counterAddrTwoStream_ready = (! counterAddrTwoStream_rValid);
  assign counterAddrTwoStream_s2mPipe_valid = (counterAddrTwoStream_valid || counterAddrTwoStream_rValid);
  assign counterAddrTwoStream_s2mPipe_payload = (counterAddrTwoStream_rValid ? counterAddrTwoStream_rData : counterAddrTwoStream_payload);
  always @(*) begin
    counterAddrTwoStream_s2mPipe_ready = counterAddrTwoStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_7) begin
      counterAddrTwoStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_7 = (! counterAddrTwoStream_s2mPipe_m2sPipe_valid);
  assign counterAddrTwoStream_s2mPipe_m2sPipe_valid = counterAddrTwoStream_s2mPipe_rValid;
  assign counterAddrTwoStream_s2mPipe_m2sPipe_payload = counterAddrTwoStream_s2mPipe_rData;
  assign counterAddrTwoStream_s2mPipe_m2sPipe_ready = ((! CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready) || CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready = CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_counterTwoPixelStream_payload = CICC1851_lineBufferTwo_port2;
  assign CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_4 = readStage_counterTwoPixelStream_ready;
    if(when_Stream_l368_8) begin
      CICC1851_4 = 1'b1;
    end
  end

  assign when_Stream_l368_8 = (! readStage_counterTwoPixelStream_valid);
  assign readStage_counterTwoPixelStream_valid = CICC1851_readStage_counterTwoPixelStream_valid;
  assign readStage_counterTwoPixelStream_payload = CICC1851_readStage_counterTwoPixelStream_payload_2;
  assign oddAddrStream_ready = (! oddAddrStream_rValid);
  assign oddAddrStream_s2mPipe_valid = (oddAddrStream_valid || oddAddrStream_rValid);
  assign oddAddrStream_s2mPipe_payload = (oddAddrStream_rValid ? oddAddrStream_rData : oddAddrStream_payload);
  always @(*) begin
    oddAddrStream_s2mPipe_ready = oddAddrStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_9) begin
      oddAddrStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_9 = (! oddAddrStream_s2mPipe_m2sPipe_valid);
  assign oddAddrStream_s2mPipe_m2sPipe_valid = oddAddrStream_s2mPipe_rValid;
  assign oddAddrStream_s2mPipe_m2sPipe_payload = oddAddrStream_s2mPipe_rData;
  assign oddAddrStream_s2mPipe_m2sPipe_ready = ((! CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready) || CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready = CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_oddRowPixelStream_payload = CICC1851_lineBufferOdd_port1;
  assign CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_5 = readStage_oddRowPixelStream_ready;
    if(when_Stream_l368_10) begin
      CICC1851_5 = 1'b1;
    end
  end

  assign when_Stream_l368_10 = (! readStage_oddRowPixelStream_valid);
  assign readStage_oddRowPixelStream_valid = CICC1851_readStage_oddRowPixelStream_valid;
  assign readStage_oddRowPixelStream_payload = CICC1851_readStage_oddRowPixelStream_payload_2;
  assign controlStream_ready = (! controlStream_rValid);
  assign controlStream_s2mPipe_valid = (controlStream_valid || controlStream_rValid);
  assign controlStream_s2mPipe_payload_frameStart = (controlStream_rValid ? controlStream_rData_frameStart : controlStream_payload_frameStart);
  assign controlStream_s2mPipe_payload_rowEnd = (controlStream_rValid ? controlStream_rData_rowEnd : controlStream_payload_rowEnd);
  assign controlStream_s2mPipe_payload_passMode = (controlStream_rValid ? controlStream_rData_passMode : controlStream_payload_passMode);
  assign controlStream_s2mPipe_payload_passValid = (controlStream_rValid ? controlStream_rData_passValid : controlStream_payload_passValid);
  assign controlStream_s2mPipe_payload_onceMode = (controlStream_rValid ? controlStream_rData_onceMode : controlStream_payload_onceMode);
  assign controlStream_s2mPipe_payload_onceValid = (controlStream_rValid ? controlStream_rData_onceValid : controlStream_payload_onceValid);
  assign controlStream_s2mPipe_payload_mainCompare = (controlStream_rValid ? controlStream_rData_mainCompare : controlStream_payload_mainCompare);
  assign controlStream_s2mPipe_payload_counterCompare = (controlStream_rValid ? controlStream_rData_counterCompare : controlStream_payload_counterCompare);
  assign controlStream_s2mPipe_payload_mainDiff = (controlStream_rValid ? controlStream_rData_mainDiff : controlStream_payload_mainDiff);
  assign controlStream_s2mPipe_payload_counterDiff = (controlStream_rValid ? controlStream_rData_counterDiff : controlStream_payload_counterDiff);
  assign controlStream_s2mPipe_payload_twiceCompValid = (controlStream_rValid ? controlStream_rData_twiceCompValid : controlStream_payload_twiceCompValid);
  assign controlStream_s2mPipe_payload_twiceMode = (controlStream_rValid ? controlStream_rData_twiceMode : controlStream_payload_twiceMode);
  assign controlStream_s2mPipe_payload_inpValidFlag = (controlStream_rValid ? controlStream_rData_inpValidFlag : controlStream_payload_inpValidFlag);
  assign controlStream_s2mPipe_payload_oddValid = (controlStream_rValid ? controlStream_rData_oddValid : controlStream_payload_oddValid);
  always @(*) begin
    controlStream_s2mPipe_ready = controlStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_11) begin
      controlStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_11 = (! controlStream_s2mPipe_m2sPipe_valid);
  assign controlStream_s2mPipe_m2sPipe_valid = controlStream_s2mPipe_rValid;
  assign controlStream_s2mPipe_m2sPipe_payload_frameStart = controlStream_s2mPipe_rData_frameStart;
  assign controlStream_s2mPipe_m2sPipe_payload_rowEnd = controlStream_s2mPipe_rData_rowEnd;
  assign controlStream_s2mPipe_m2sPipe_payload_passMode = controlStream_s2mPipe_rData_passMode;
  assign controlStream_s2mPipe_m2sPipe_payload_passValid = controlStream_s2mPipe_rData_passValid;
  assign controlStream_s2mPipe_m2sPipe_payload_onceMode = controlStream_s2mPipe_rData_onceMode;
  assign controlStream_s2mPipe_m2sPipe_payload_onceValid = controlStream_s2mPipe_rData_onceValid;
  assign controlStream_s2mPipe_m2sPipe_payload_mainCompare = controlStream_s2mPipe_rData_mainCompare;
  assign controlStream_s2mPipe_m2sPipe_payload_counterCompare = controlStream_s2mPipe_rData_counterCompare;
  assign controlStream_s2mPipe_m2sPipe_payload_mainDiff = controlStream_s2mPipe_rData_mainDiff;
  assign controlStream_s2mPipe_m2sPipe_payload_counterDiff = controlStream_s2mPipe_rData_counterDiff;
  assign controlStream_s2mPipe_m2sPipe_payload_twiceCompValid = controlStream_s2mPipe_rData_twiceCompValid;
  assign controlStream_s2mPipe_m2sPipe_payload_twiceMode = controlStream_s2mPipe_rData_twiceMode;
  assign controlStream_s2mPipe_m2sPipe_payload_inpValidFlag = controlStream_s2mPipe_rData_inpValidFlag;
  assign controlStream_s2mPipe_m2sPipe_payload_oddValid = controlStream_s2mPipe_rData_oddValid;
  always @(*) begin
    controlStream_s2mPipe_m2sPipe_ready = controlStream_s2mPipe_m2sPipe_m2sPipe_ready;
    if(when_Stream_l368_12) begin
      controlStream_s2mPipe_m2sPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_12 = (! controlStream_s2mPipe_m2sPipe_m2sPipe_valid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_valid = controlStream_s2mPipe_m2sPipe_rValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_frameStart = controlStream_s2mPipe_m2sPipe_rData_frameStart;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_rowEnd = controlStream_s2mPipe_m2sPipe_rData_rowEnd;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passMode = controlStream_s2mPipe_m2sPipe_rData_passMode;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passValid = controlStream_s2mPipe_m2sPipe_rData_passValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceMode = controlStream_s2mPipe_m2sPipe_rData_onceMode;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceValid = controlStream_s2mPipe_m2sPipe_rData_onceValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainCompare = controlStream_s2mPipe_m2sPipe_rData_mainCompare;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterCompare = controlStream_s2mPipe_m2sPipe_rData_counterCompare;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDiff = controlStream_s2mPipe_m2sPipe_rData_mainDiff;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDiff = controlStream_s2mPipe_m2sPipe_rData_counterDiff;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceCompValid = controlStream_s2mPipe_m2sPipe_rData_twiceCompValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceMode = controlStream_s2mPipe_m2sPipe_rData_twiceMode;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_inpValidFlag = controlStream_s2mPipe_m2sPipe_rData_inpValidFlag;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_oddValid = controlStream_s2mPipe_m2sPipe_rData_oddValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_ready = (! controlStream_s2mPipe_m2sPipe_m2sPipe_rValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_valid = (controlStream_s2mPipe_m2sPipe_m2sPipe_valid || controlStream_s2mPipe_m2sPipe_m2sPipe_rValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_frameStart = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_frameStart : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_frameStart);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_rowEnd = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_rowEnd : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_rowEnd);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_passMode = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_passMode : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passMode);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_passValid = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_passValid : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_onceMode = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_onceMode : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceMode);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_onceValid = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_onceValid : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainCompare = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainCompare : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainCompare);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterCompare = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterCompare : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterCompare);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainDiff = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainDiff : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDiff);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterDiff = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterDiff : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDiff);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_twiceCompValid = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_twiceCompValid : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceCompValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_twiceMode = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_twiceMode : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceMode);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_inpValidFlag = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_inpValidFlag : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_inpValidFlag);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_oddValid = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_oddValid : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_oddValid);
  always @(*) begin
    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready = readStage_controlPipe_ready;
    if(when_Stream_l368_13) begin
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_13 = (! readStage_controlPipe_valid);
  assign readStage_controlPipe_valid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rValid;
  assign readStage_controlPipe_payload_frameStart = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_frameStart;
  assign readStage_controlPipe_payload_rowEnd = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_rowEnd;
  assign readStage_controlPipe_payload_passMode = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_passMode;
  assign readStage_controlPipe_payload_passValid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_passValid;
  assign readStage_controlPipe_payload_onceMode = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_onceMode;
  assign readStage_controlPipe_payload_onceValid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_onceValid;
  assign readStage_controlPipe_payload_mainCompare = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainCompare;
  assign readStage_controlPipe_payload_counterCompare = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterCompare;
  assign readStage_controlPipe_payload_mainDiff = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainDiff;
  assign readStage_controlPipe_payload_counterDiff = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterDiff;
  assign readStage_controlPipe_payload_twiceCompValid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_twiceCompValid;
  assign readStage_controlPipe_payload_twiceMode = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_twiceMode;
  assign readStage_controlPipe_payload_inpValidFlag = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_inpValidFlag;
  assign readStage_controlPipe_payload_oddValid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_oddValid;
  assign readStage_mainOnePixelStream_ready = (! readStage_mainOnePixelStream_rValid);
  assign readStage_mainOnePixelStream_s2mPipe_valid = (readStage_mainOnePixelStream_valid || readStage_mainOnePixelStream_rValid);
  assign readStage_mainOnePixelStream_s2mPipe_payload = (readStage_mainOnePixelStream_rValid ? readStage_mainOnePixelStream_rData : readStage_mainOnePixelStream_payload);
  always @(*) begin
    readStage_mainOnePixelStream_s2mPipe_ready = compareStage_mainOnePixelStream_ready;
    if(when_Stream_l368_14) begin
      readStage_mainOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_14 = (! compareStage_mainOnePixelStream_valid);
  assign compareStage_mainOnePixelStream_valid = readStage_mainOnePixelStream_s2mPipe_rValid;
  assign compareStage_mainOnePixelStream_payload = readStage_mainOnePixelStream_s2mPipe_rData;
  assign readStage_counterOnePixelStream_ready = (! readStage_counterOnePixelStream_rValid);
  assign readStage_counterOnePixelStream_s2mPipe_valid = (readStage_counterOnePixelStream_valid || readStage_counterOnePixelStream_rValid);
  assign readStage_counterOnePixelStream_s2mPipe_payload = (readStage_counterOnePixelStream_rValid ? readStage_counterOnePixelStream_rData : readStage_counterOnePixelStream_payload);
  always @(*) begin
    readStage_counterOnePixelStream_s2mPipe_ready = compareStage_counterOnePixelStream_ready;
    if(when_Stream_l368_15) begin
      readStage_counterOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_15 = (! compareStage_counterOnePixelStream_valid);
  assign compareStage_counterOnePixelStream_valid = readStage_counterOnePixelStream_s2mPipe_rValid;
  assign compareStage_counterOnePixelStream_payload = readStage_counterOnePixelStream_s2mPipe_rData;
  assign readStage_mainTwoPixelStream_ready = (! readStage_mainTwoPixelStream_rValid);
  assign readStage_mainTwoPixelStream_s2mPipe_valid = (readStage_mainTwoPixelStream_valid || readStage_mainTwoPixelStream_rValid);
  assign readStage_mainTwoPixelStream_s2mPipe_payload = (readStage_mainTwoPixelStream_rValid ? readStage_mainTwoPixelStream_rData : readStage_mainTwoPixelStream_payload);
  always @(*) begin
    readStage_mainTwoPixelStream_s2mPipe_ready = compareStage_mainTwoPixelStream_ready;
    if(when_Stream_l368_16) begin
      readStage_mainTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_16 = (! compareStage_mainTwoPixelStream_valid);
  assign compareStage_mainTwoPixelStream_valid = readStage_mainTwoPixelStream_s2mPipe_rValid;
  assign compareStage_mainTwoPixelStream_payload = readStage_mainTwoPixelStream_s2mPipe_rData;
  assign readStage_counterTwoPixelStream_ready = (! readStage_counterTwoPixelStream_rValid);
  assign readStage_counterTwoPixelStream_s2mPipe_valid = (readStage_counterTwoPixelStream_valid || readStage_counterTwoPixelStream_rValid);
  assign readStage_counterTwoPixelStream_s2mPipe_payload = (readStage_counterTwoPixelStream_rValid ? readStage_counterTwoPixelStream_rData : readStage_counterTwoPixelStream_payload);
  always @(*) begin
    readStage_counterTwoPixelStream_s2mPipe_ready = compareStage_counterTwoPixelStream_ready;
    if(when_Stream_l368_17) begin
      readStage_counterTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_17 = (! compareStage_counterTwoPixelStream_valid);
  assign compareStage_counterTwoPixelStream_valid = readStage_counterTwoPixelStream_s2mPipe_rValid;
  assign compareStage_counterTwoPixelStream_payload = readStage_counterTwoPixelStream_s2mPipe_rData;
  assign readStage_oddRowPixelStream_ready = (! readStage_oddRowPixelStream_rValid);
  assign readStage_oddRowPixelStream_s2mPipe_valid = (readStage_oddRowPixelStream_valid || readStage_oddRowPixelStream_rValid);
  assign readStage_oddRowPixelStream_s2mPipe_payload = (readStage_oddRowPixelStream_rValid ? readStage_oddRowPixelStream_rData : readStage_oddRowPixelStream_payload);
  always @(*) begin
    readStage_oddRowPixelStream_s2mPipe_ready = compareStage_oddRowPixelStream_ready;
    if(when_Stream_l368_18) begin
      readStage_oddRowPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_18 = (! compareStage_oddRowPixelStream_valid);
  assign compareStage_oddRowPixelStream_valid = readStage_oddRowPixelStream_s2mPipe_rValid;
  assign compareStage_oddRowPixelStream_payload = readStage_oddRowPixelStream_s2mPipe_rData;
  always @(*) begin
    CICC1851_readStage_controlPipe_translated_payload_mainCompare = readStage_controlPipe_payload_mainCompare;
    if(readStage_controlPipe_payload_onceValid) begin
      case(readStage_controlPipe_payload_onceMode)
        3'b000 : begin
          if(when_SuperResolutionPart2_l290) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        3'b001 : begin
          if(when_SuperResolutionPart2_l294) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        3'b010 : begin
          if(when_SuperResolutionPart2_l298) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        3'b011 : begin
          if(when_SuperResolutionPart2_l302) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        3'b100 : begin
          CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
        end
        3'b101 : begin
          CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
        end
        default : begin
        end
      endcase
    end
    if(readStage_controlPipe_payload_twiceCompValid) begin
      case(readStage_controlPipe_payload_twiceMode)
        3'b000 : begin
          if(when_SuperResolutionPart2_l313) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        3'b001 : begin
          if(when_SuperResolutionPart2_l319) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        3'b010 : begin
          CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
        end
        3'b011 : begin
          if(when_SuperResolutionPart2_l326) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        3'b100 : begin
          CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
        end
        3'b101 : begin
          if(when_SuperResolutionPart2_l331) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    CICC1851_readStage_controlPipe_translated_payload_counterCompare = readStage_controlPipe_payload_counterCompare;
    if(readStage_controlPipe_payload_twiceCompValid) begin
      case(readStage_controlPipe_payload_twiceMode)
        3'b000 : begin
          if(when_SuperResolutionPart2_l315) begin
            CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
          end
        end
        3'b001 : begin
          if(when_SuperResolutionPart2_l321) begin
            CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
          end
        end
        default : begin
        end
      endcase
    end
  end

  assign when_SuperResolutionPart2_l290 = (readStage_counterOnePixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart2_l294 = (readStage_counterTwoPixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart2_l298 = (readStage_mainTwoPixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart2_l302 = (readStage_mainOnePixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart2_l313 = (readStage_mainTwoPixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart2_l315 = (readStage_counterOnePixelStream_payload <= readStage_counterTwoPixelStream_payload);
  assign when_SuperResolutionPart2_l319 = (readStage_mainOnePixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart2_l321 = (readStage_counterTwoPixelStream_payload <= readStage_counterOnePixelStream_payload);
  assign when_SuperResolutionPart2_l326 = (readStage_counterTwoPixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart2_l331 = (readStage_counterOnePixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign readStage_controlPipe_translated_valid = readStage_controlPipe_valid;
  assign readStage_controlPipe_ready = readStage_controlPipe_translated_ready;
  assign readStage_controlPipe_translated_payload_frameStart = readStage_controlPipe_payload_frameStart;
  assign readStage_controlPipe_translated_payload_rowEnd = readStage_controlPipe_payload_rowEnd;
  assign readStage_controlPipe_translated_payload_passMode = readStage_controlPipe_payload_passMode;
  assign readStage_controlPipe_translated_payload_passValid = readStage_controlPipe_payload_passValid;
  assign readStage_controlPipe_translated_payload_onceMode = readStage_controlPipe_payload_onceMode;
  assign readStage_controlPipe_translated_payload_onceValid = readStage_controlPipe_payload_onceValid;
  assign readStage_controlPipe_translated_payload_mainCompare = CICC1851_readStage_controlPipe_translated_payload_mainCompare;
  assign readStage_controlPipe_translated_payload_counterCompare = CICC1851_readStage_controlPipe_translated_payload_counterCompare;
  assign readStage_controlPipe_translated_payload_mainDiff = readStage_controlPipe_payload_mainDiff;
  assign readStage_controlPipe_translated_payload_counterDiff = readStage_controlPipe_payload_counterDiff;
  assign readStage_controlPipe_translated_payload_twiceCompValid = readStage_controlPipe_payload_twiceCompValid;
  assign readStage_controlPipe_translated_payload_twiceMode = readStage_controlPipe_payload_twiceMode;
  assign readStage_controlPipe_translated_payload_inpValidFlag = readStage_controlPipe_payload_inpValidFlag;
  assign readStage_controlPipe_translated_payload_oddValid = readStage_controlPipe_payload_oddValid;
  assign readStage_controlPipe_translated_ready = (! readStage_controlPipe_translated_rValid);
  assign readStage_controlPipe_translated_s2mPipe_valid = (readStage_controlPipe_translated_valid || readStage_controlPipe_translated_rValid);
  assign readStage_controlPipe_translated_s2mPipe_payload_frameStart = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_frameStart : readStage_controlPipe_translated_payload_frameStart);
  assign readStage_controlPipe_translated_s2mPipe_payload_rowEnd = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_rowEnd : readStage_controlPipe_translated_payload_rowEnd);
  assign readStage_controlPipe_translated_s2mPipe_payload_passMode = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_passMode : readStage_controlPipe_translated_payload_passMode);
  assign readStage_controlPipe_translated_s2mPipe_payload_passValid = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_passValid : readStage_controlPipe_translated_payload_passValid);
  assign readStage_controlPipe_translated_s2mPipe_payload_onceMode = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_onceMode : readStage_controlPipe_translated_payload_onceMode);
  assign readStage_controlPipe_translated_s2mPipe_payload_onceValid = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_onceValid : readStage_controlPipe_translated_payload_onceValid);
  assign readStage_controlPipe_translated_s2mPipe_payload_mainCompare = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_mainCompare : readStage_controlPipe_translated_payload_mainCompare);
  assign readStage_controlPipe_translated_s2mPipe_payload_counterCompare = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_counterCompare : readStage_controlPipe_translated_payload_counterCompare);
  assign readStage_controlPipe_translated_s2mPipe_payload_mainDiff = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_mainDiff : readStage_controlPipe_translated_payload_mainDiff);
  assign readStage_controlPipe_translated_s2mPipe_payload_counterDiff = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_counterDiff : readStage_controlPipe_translated_payload_counterDiff);
  assign readStage_controlPipe_translated_s2mPipe_payload_twiceCompValid = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_twiceCompValid : readStage_controlPipe_translated_payload_twiceCompValid);
  assign readStage_controlPipe_translated_s2mPipe_payload_twiceMode = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_twiceMode : readStage_controlPipe_translated_payload_twiceMode);
  assign readStage_controlPipe_translated_s2mPipe_payload_inpValidFlag = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_inpValidFlag : readStage_controlPipe_translated_payload_inpValidFlag);
  assign readStage_controlPipe_translated_s2mPipe_payload_oddValid = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_oddValid : readStage_controlPipe_translated_payload_oddValid);
  always @(*) begin
    readStage_controlPipe_translated_s2mPipe_ready = compareStage_controlPipe_ready;
    if(when_Stream_l368_19) begin
      readStage_controlPipe_translated_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_19 = (! compareStage_controlPipe_valid);
  assign compareStage_controlPipe_valid = readStage_controlPipe_translated_s2mPipe_rValid;
  assign compareStage_controlPipe_payload_frameStart = readStage_controlPipe_translated_s2mPipe_rData_frameStart;
  assign compareStage_controlPipe_payload_rowEnd = readStage_controlPipe_translated_s2mPipe_rData_rowEnd;
  assign compareStage_controlPipe_payload_passMode = readStage_controlPipe_translated_s2mPipe_rData_passMode;
  assign compareStage_controlPipe_payload_passValid = readStage_controlPipe_translated_s2mPipe_rData_passValid;
  assign compareStage_controlPipe_payload_onceMode = readStage_controlPipe_translated_s2mPipe_rData_onceMode;
  assign compareStage_controlPipe_payload_onceValid = readStage_controlPipe_translated_s2mPipe_rData_onceValid;
  assign compareStage_controlPipe_payload_mainCompare = readStage_controlPipe_translated_s2mPipe_rData_mainCompare;
  assign compareStage_controlPipe_payload_counterCompare = readStage_controlPipe_translated_s2mPipe_rData_counterCompare;
  assign compareStage_controlPipe_payload_mainDiff = readStage_controlPipe_translated_s2mPipe_rData_mainDiff;
  assign compareStage_controlPipe_payload_counterDiff = readStage_controlPipe_translated_s2mPipe_rData_counterDiff;
  assign compareStage_controlPipe_payload_twiceCompValid = readStage_controlPipe_translated_s2mPipe_rData_twiceCompValid;
  assign compareStage_controlPipe_payload_twiceMode = readStage_controlPipe_translated_s2mPipe_rData_twiceMode;
  assign compareStage_controlPipe_payload_inpValidFlag = readStage_controlPipe_translated_s2mPipe_rData_inpValidFlag;
  assign compareStage_controlPipe_payload_oddValid = readStage_controlPipe_translated_s2mPipe_rData_oddValid;
  assign compareStage_mainOnePixelStream_ready = (! compareStage_mainOnePixelStream_rValid);
  assign compareStage_mainOnePixelStream_s2mPipe_valid = (compareStage_mainOnePixelStream_valid || compareStage_mainOnePixelStream_rValid);
  assign compareStage_mainOnePixelStream_s2mPipe_payload = (compareStage_mainOnePixelStream_rValid ? compareStage_mainOnePixelStream_rData : compareStage_mainOnePixelStream_payload);
  always @(*) begin
    compareStage_mainOnePixelStream_s2mPipe_ready = diffStage_mainOnePixelStream_ready;
    if(when_Stream_l368_20) begin
      compareStage_mainOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_20 = (! diffStage_mainOnePixelStream_valid);
  assign diffStage_mainOnePixelStream_valid = compareStage_mainOnePixelStream_s2mPipe_rValid;
  assign diffStage_mainOnePixelStream_payload = compareStage_mainOnePixelStream_s2mPipe_rData;
  assign compareStage_counterOnePixelStream_ready = (! compareStage_counterOnePixelStream_rValid);
  assign compareStage_counterOnePixelStream_s2mPipe_valid = (compareStage_counterOnePixelStream_valid || compareStage_counterOnePixelStream_rValid);
  assign compareStage_counterOnePixelStream_s2mPipe_payload = (compareStage_counterOnePixelStream_rValid ? compareStage_counterOnePixelStream_rData : compareStage_counterOnePixelStream_payload);
  always @(*) begin
    compareStage_counterOnePixelStream_s2mPipe_ready = diffStage_counterOnePixelStream_ready;
    if(when_Stream_l368_21) begin
      compareStage_counterOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_21 = (! diffStage_counterOnePixelStream_valid);
  assign diffStage_counterOnePixelStream_valid = compareStage_counterOnePixelStream_s2mPipe_rValid;
  assign diffStage_counterOnePixelStream_payload = compareStage_counterOnePixelStream_s2mPipe_rData;
  assign compareStage_mainTwoPixelStream_ready = (! compareStage_mainTwoPixelStream_rValid);
  assign compareStage_mainTwoPixelStream_s2mPipe_valid = (compareStage_mainTwoPixelStream_valid || compareStage_mainTwoPixelStream_rValid);
  assign compareStage_mainTwoPixelStream_s2mPipe_payload = (compareStage_mainTwoPixelStream_rValid ? compareStage_mainTwoPixelStream_rData : compareStage_mainTwoPixelStream_payload);
  always @(*) begin
    compareStage_mainTwoPixelStream_s2mPipe_ready = diffStage_mainTwoPixelStream_ready;
    if(when_Stream_l368_22) begin
      compareStage_mainTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_22 = (! diffStage_mainTwoPixelStream_valid);
  assign diffStage_mainTwoPixelStream_valid = compareStage_mainTwoPixelStream_s2mPipe_rValid;
  assign diffStage_mainTwoPixelStream_payload = compareStage_mainTwoPixelStream_s2mPipe_rData;
  assign compareStage_counterTwoPixelStream_ready = (! compareStage_counterTwoPixelStream_rValid);
  assign compareStage_counterTwoPixelStream_s2mPipe_valid = (compareStage_counterTwoPixelStream_valid || compareStage_counterTwoPixelStream_rValid);
  assign compareStage_counterTwoPixelStream_s2mPipe_payload = (compareStage_counterTwoPixelStream_rValid ? compareStage_counterTwoPixelStream_rData : compareStage_counterTwoPixelStream_payload);
  always @(*) begin
    compareStage_counterTwoPixelStream_s2mPipe_ready = diffStage_counterTwoPixelStream_ready;
    if(when_Stream_l368_23) begin
      compareStage_counterTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_23 = (! diffStage_counterTwoPixelStream_valid);
  assign diffStage_counterTwoPixelStream_valid = compareStage_counterTwoPixelStream_s2mPipe_rValid;
  assign diffStage_counterTwoPixelStream_payload = compareStage_counterTwoPixelStream_s2mPipe_rData;
  assign compareStage_oddRowPixelStream_ready = (! compareStage_oddRowPixelStream_rValid);
  assign compareStage_oddRowPixelStream_s2mPipe_valid = (compareStage_oddRowPixelStream_valid || compareStage_oddRowPixelStream_rValid);
  assign compareStage_oddRowPixelStream_s2mPipe_payload = (compareStage_oddRowPixelStream_rValid ? compareStage_oddRowPixelStream_rData : compareStage_oddRowPixelStream_payload);
  always @(*) begin
    compareStage_oddRowPixelStream_s2mPipe_ready = diffStage_oddRowPixelStream_ready;
    if(when_Stream_l368_24) begin
      compareStage_oddRowPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_24 = (! diffStage_oddRowPixelStream_valid);
  assign diffStage_oddRowPixelStream_valid = compareStage_oddRowPixelStream_s2mPipe_rValid;
  assign diffStage_oddRowPixelStream_payload = compareStage_oddRowPixelStream_s2mPipe_rData;
  always @(*) begin
    CICC1851_compareStage_controlPipe_translated_payload_mainDiff = compareStage_controlPipe_payload_mainDiff;
    if(compareStage_controlPipe_payload_onceValid) begin
      case(compareStage_controlPipe_payload_onceMode)
        3'b000 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_counterOnePixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterOnePixelStream_payload - compareStage_mainOnePixelStream_payload);
          end
        end
        3'b001 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterTwoPixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainTwoPixelStream_payload);
          end
        end
        3'b010 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_mainTwoPixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_mainOnePixelStream_payload);
          end
        end
        3'b011 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_mainOnePixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_mainTwoPixelStream_payload);
          end
        end
        3'b100 : begin
          CICC1851_compareStage_controlPipe_translated_payload_mainDiff = 8'h0;
        end
        3'b101 : begin
          CICC1851_compareStage_controlPipe_translated_payload_mainDiff = 8'h0;
        end
        default : begin
        end
      endcase
    end
    if(compareStage_controlPipe_payload_twiceCompValid) begin
      case(compareStage_controlPipe_payload_twiceMode)
        3'b000 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_mainTwoPixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_mainOnePixelStream_payload);
          end
        end
        3'b001 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_mainOnePixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_mainTwoPixelStream_payload);
          end
        end
        3'b010 : begin
          CICC1851_compareStage_controlPipe_translated_payload_mainDiff = 8'h0;
        end
        3'b011 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterTwoPixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainTwoPixelStream_payload);
          end
        end
        3'b100 : begin
          CICC1851_compareStage_controlPipe_translated_payload_mainDiff = 8'h0;
        end
        3'b101 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_counterOnePixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterOnePixelStream_payload - compareStage_mainOnePixelStream_payload);
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    CICC1851_compareStage_controlPipe_translated_payload_counterDiff = compareStage_controlPipe_payload_counterDiff;
    if(compareStage_controlPipe_payload_twiceCompValid) begin
      case(compareStage_controlPipe_payload_twiceMode)
        3'b000 : begin
          if(compareStage_controlPipe_payload_counterCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterTwoPixelStream_payload - compareStage_counterOnePixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterOnePixelStream_payload - compareStage_counterTwoPixelStream_payload);
          end
        end
        3'b001 : begin
          if(compareStage_controlPipe_payload_counterCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterOnePixelStream_payload - compareStage_counterTwoPixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterTwoPixelStream_payload - compareStage_counterOnePixelStream_payload);
          end
        end
        default : begin
        end
      endcase
    end
  end

  assign compareStage_controlPipe_translated_valid = compareStage_controlPipe_valid;
  assign compareStage_controlPipe_ready = compareStage_controlPipe_translated_ready;
  assign compareStage_controlPipe_translated_payload_frameStart = compareStage_controlPipe_payload_frameStart;
  assign compareStage_controlPipe_translated_payload_rowEnd = compareStage_controlPipe_payload_rowEnd;
  assign compareStage_controlPipe_translated_payload_passMode = compareStage_controlPipe_payload_passMode;
  assign compareStage_controlPipe_translated_payload_passValid = compareStage_controlPipe_payload_passValid;
  assign compareStage_controlPipe_translated_payload_onceMode = compareStage_controlPipe_payload_onceMode;
  assign compareStage_controlPipe_translated_payload_onceValid = compareStage_controlPipe_payload_onceValid;
  assign compareStage_controlPipe_translated_payload_mainCompare = compareStage_controlPipe_payload_mainCompare;
  assign compareStage_controlPipe_translated_payload_counterCompare = compareStage_controlPipe_payload_counterCompare;
  assign compareStage_controlPipe_translated_payload_mainDiff = CICC1851_compareStage_controlPipe_translated_payload_mainDiff;
  assign compareStage_controlPipe_translated_payload_counterDiff = CICC1851_compareStage_controlPipe_translated_payload_counterDiff;
  assign compareStage_controlPipe_translated_payload_twiceCompValid = compareStage_controlPipe_payload_twiceCompValid;
  assign compareStage_controlPipe_translated_payload_twiceMode = compareStage_controlPipe_payload_twiceMode;
  assign compareStage_controlPipe_translated_payload_inpValidFlag = compareStage_controlPipe_payload_inpValidFlag;
  assign compareStage_controlPipe_translated_payload_oddValid = compareStage_controlPipe_payload_oddValid;
  assign compareStage_controlPipe_translated_ready = (! compareStage_controlPipe_translated_rValid);
  assign compareStage_controlPipe_translated_s2mPipe_valid = (compareStage_controlPipe_translated_valid || compareStage_controlPipe_translated_rValid);
  assign compareStage_controlPipe_translated_s2mPipe_payload_frameStart = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_frameStart : compareStage_controlPipe_translated_payload_frameStart);
  assign compareStage_controlPipe_translated_s2mPipe_payload_rowEnd = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_rowEnd : compareStage_controlPipe_translated_payload_rowEnd);
  assign compareStage_controlPipe_translated_s2mPipe_payload_passMode = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_passMode : compareStage_controlPipe_translated_payload_passMode);
  assign compareStage_controlPipe_translated_s2mPipe_payload_passValid = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_passValid : compareStage_controlPipe_translated_payload_passValid);
  assign compareStage_controlPipe_translated_s2mPipe_payload_onceMode = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_onceMode : compareStage_controlPipe_translated_payload_onceMode);
  assign compareStage_controlPipe_translated_s2mPipe_payload_onceValid = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_onceValid : compareStage_controlPipe_translated_payload_onceValid);
  assign compareStage_controlPipe_translated_s2mPipe_payload_mainCompare = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_mainCompare : compareStage_controlPipe_translated_payload_mainCompare);
  assign compareStage_controlPipe_translated_s2mPipe_payload_counterCompare = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_counterCompare : compareStage_controlPipe_translated_payload_counterCompare);
  assign compareStage_controlPipe_translated_s2mPipe_payload_mainDiff = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_mainDiff : compareStage_controlPipe_translated_payload_mainDiff);
  assign compareStage_controlPipe_translated_s2mPipe_payload_counterDiff = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_counterDiff : compareStage_controlPipe_translated_payload_counterDiff);
  assign compareStage_controlPipe_translated_s2mPipe_payload_twiceCompValid = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_twiceCompValid : compareStage_controlPipe_translated_payload_twiceCompValid);
  assign compareStage_controlPipe_translated_s2mPipe_payload_twiceMode = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_twiceMode : compareStage_controlPipe_translated_payload_twiceMode);
  assign compareStage_controlPipe_translated_s2mPipe_payload_inpValidFlag = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_inpValidFlag : compareStage_controlPipe_translated_payload_inpValidFlag);
  assign compareStage_controlPipe_translated_s2mPipe_payload_oddValid = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_oddValid : compareStage_controlPipe_translated_payload_oddValid);
  always @(*) begin
    compareStage_controlPipe_translated_s2mPipe_ready = diffStage_controlPipe_ready;
    if(when_Stream_l368_25) begin
      compareStage_controlPipe_translated_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_25 = (! diffStage_controlPipe_valid);
  assign diffStage_controlPipe_valid = compareStage_controlPipe_translated_s2mPipe_rValid;
  assign diffStage_controlPipe_payload_frameStart = compareStage_controlPipe_translated_s2mPipe_rData_frameStart;
  assign diffStage_controlPipe_payload_rowEnd = compareStage_controlPipe_translated_s2mPipe_rData_rowEnd;
  assign diffStage_controlPipe_payload_passMode = compareStage_controlPipe_translated_s2mPipe_rData_passMode;
  assign diffStage_controlPipe_payload_passValid = compareStage_controlPipe_translated_s2mPipe_rData_passValid;
  assign diffStage_controlPipe_payload_onceMode = compareStage_controlPipe_translated_s2mPipe_rData_onceMode;
  assign diffStage_controlPipe_payload_onceValid = compareStage_controlPipe_translated_s2mPipe_rData_onceValid;
  assign diffStage_controlPipe_payload_mainCompare = compareStage_controlPipe_translated_s2mPipe_rData_mainCompare;
  assign diffStage_controlPipe_payload_counterCompare = compareStage_controlPipe_translated_s2mPipe_rData_counterCompare;
  assign diffStage_controlPipe_payload_mainDiff = compareStage_controlPipe_translated_s2mPipe_rData_mainDiff;
  assign diffStage_controlPipe_payload_counterDiff = compareStage_controlPipe_translated_s2mPipe_rData_counterDiff;
  assign diffStage_controlPipe_payload_twiceCompValid = compareStage_controlPipe_translated_s2mPipe_rData_twiceCompValid;
  assign diffStage_controlPipe_payload_twiceMode = compareStage_controlPipe_translated_s2mPipe_rData_twiceMode;
  assign diffStage_controlPipe_payload_inpValidFlag = compareStage_controlPipe_translated_s2mPipe_rData_inpValidFlag;
  assign diffStage_controlPipe_payload_oddValid = compareStage_controlPipe_translated_s2mPipe_rData_oddValid;
  assign diffStage_mainOnePixelStream_ready = (! diffStage_mainOnePixelStream_rValid);
  assign diffStage_mainOnePixelStream_s2mPipe_valid = (diffStage_mainOnePixelStream_valid || diffStage_mainOnePixelStream_rValid);
  assign diffStage_mainOnePixelStream_s2mPipe_payload = (diffStage_mainOnePixelStream_rValid ? diffStage_mainOnePixelStream_rData : diffStage_mainOnePixelStream_payload);
  always @(*) begin
    diffStage_mainOnePixelStream_s2mPipe_ready = resultStage_mainOnePixelStream_ready;
    if(when_Stream_l368_26) begin
      diffStage_mainOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_26 = (! resultStage_mainOnePixelStream_valid);
  assign resultStage_mainOnePixelStream_valid = diffStage_mainOnePixelStream_s2mPipe_rValid;
  assign resultStage_mainOnePixelStream_payload = diffStage_mainOnePixelStream_s2mPipe_rData;
  assign diffStage_counterOnePixelStream_ready = (! diffStage_counterOnePixelStream_rValid);
  assign diffStage_counterOnePixelStream_s2mPipe_valid = (diffStage_counterOnePixelStream_valid || diffStage_counterOnePixelStream_rValid);
  assign diffStage_counterOnePixelStream_s2mPipe_payload = (diffStage_counterOnePixelStream_rValid ? diffStage_counterOnePixelStream_rData : diffStage_counterOnePixelStream_payload);
  always @(*) begin
    diffStage_counterOnePixelStream_s2mPipe_ready = resultStage_counterOnePixelStream_ready;
    if(when_Stream_l368_27) begin
      diffStage_counterOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_27 = (! resultStage_counterOnePixelStream_valid);
  assign resultStage_counterOnePixelStream_valid = diffStage_counterOnePixelStream_s2mPipe_rValid;
  assign resultStage_counterOnePixelStream_payload = diffStage_counterOnePixelStream_s2mPipe_rData;
  assign diffStage_mainTwoPixelStream_ready = (! diffStage_mainTwoPixelStream_rValid);
  assign diffStage_mainTwoPixelStream_s2mPipe_valid = (diffStage_mainTwoPixelStream_valid || diffStage_mainTwoPixelStream_rValid);
  assign diffStage_mainTwoPixelStream_s2mPipe_payload = (diffStage_mainTwoPixelStream_rValid ? diffStage_mainTwoPixelStream_rData : diffStage_mainTwoPixelStream_payload);
  always @(*) begin
    diffStage_mainTwoPixelStream_s2mPipe_ready = resultStage_mainTwoPixelStream_ready;
    if(when_Stream_l368_28) begin
      diffStage_mainTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_28 = (! resultStage_mainTwoPixelStream_valid);
  assign resultStage_mainTwoPixelStream_valid = diffStage_mainTwoPixelStream_s2mPipe_rValid;
  assign resultStage_mainTwoPixelStream_payload = diffStage_mainTwoPixelStream_s2mPipe_rData;
  assign diffStage_counterTwoPixelStream_ready = (! diffStage_counterTwoPixelStream_rValid);
  assign diffStage_counterTwoPixelStream_s2mPipe_valid = (diffStage_counterTwoPixelStream_valid || diffStage_counterTwoPixelStream_rValid);
  assign diffStage_counterTwoPixelStream_s2mPipe_payload = (diffStage_counterTwoPixelStream_rValid ? diffStage_counterTwoPixelStream_rData : diffStage_counterTwoPixelStream_payload);
  always @(*) begin
    diffStage_counterTwoPixelStream_s2mPipe_ready = resultStage_counterTwoPixelStream_ready;
    if(when_Stream_l368_29) begin
      diffStage_counterTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_29 = (! resultStage_counterTwoPixelStream_valid);
  assign resultStage_counterTwoPixelStream_valid = diffStage_counterTwoPixelStream_s2mPipe_rValid;
  assign resultStage_counterTwoPixelStream_payload = diffStage_counterTwoPixelStream_s2mPipe_rData;
  assign diffStage_oddRowPixelStream_ready = (! diffStage_oddRowPixelStream_rValid);
  assign diffStage_oddRowPixelStream_s2mPipe_valid = (diffStage_oddRowPixelStream_valid || diffStage_oddRowPixelStream_rValid);
  assign diffStage_oddRowPixelStream_s2mPipe_payload = (diffStage_oddRowPixelStream_rValid ? diffStage_oddRowPixelStream_rData : diffStage_oddRowPixelStream_payload);
  always @(*) begin
    diffStage_oddRowPixelStream_s2mPipe_ready = resultStage_oddRowPixelStream_ready;
    if(when_Stream_l368_30) begin
      diffStage_oddRowPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_30 = (! resultStage_oddRowPixelStream_valid);
  assign resultStage_oddRowPixelStream_valid = diffStage_oddRowPixelStream_s2mPipe_rValid;
  assign resultStage_oddRowPixelStream_payload = diffStage_oddRowPixelStream_s2mPipe_rData;
  assign diffStage_controlPipe_ready = diffStage_controlPipe_fork_io_input_ready;
  assign CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceMode = diffStage_controlPipe_payload_onceMode;
  assign CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceValid = diffStage_controlPipe_payload_onceValid;
  assign CICC1851_when_SuperResolutionPart2_l419 = diffStage_controlPipe_payload_mainDiff;
  assign CICC1851_when_SuperResolutionPart2_l428 = diffStage_controlPipe_payload_counterDiff;
  assign CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceCompValid = diffStage_controlPipe_payload_twiceCompValid;
  assign CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceMode = diffStage_controlPipe_payload_twiceMode;
  always @(*) begin
    CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag = diffStage_controlPipe_payload_inpValidFlag;
    if(CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceValid) begin
      case(CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceMode)
        3'b000 : begin
          if(when_SuperResolutionPart2_l419) begin
            CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag = 1'b0;
          end
        end
        3'b001 : begin
          if(when_SuperResolutionPart2_l420) begin
            CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag = 1'b0;
          end
        end
        3'b010 : begin
          if(when_SuperResolutionPart2_l421) begin
            CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag = 1'b0;
          end
        end
        3'b011 : begin
          if(when_SuperResolutionPart2_l422) begin
            CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag = 1'b0;
          end
        end
        default : begin
        end
      endcase
    end
    if(CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceCompValid) begin
      case(CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceMode)
        3'b000 : begin
          if(when_SuperResolutionPart2_l428) begin
            CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag = 1'b0;
          end
        end
        3'b001 : begin
          if(when_SuperResolutionPart2_l429) begin
            CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag = 1'b0;
          end
        end
        3'b011 : begin
          if(when_SuperResolutionPart2_l430) begin
            CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag = 1'b0;
          end
        end
        3'b101 : begin
          if(when_SuperResolutionPart2_l431) begin
            CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag = 1'b0;
          end
        end
        default : begin
        end
      endcase
    end
  end

  assign when_SuperResolutionPart2_l419 = (inpThreshold <= CICC1851_when_SuperResolutionPart2_l419);
  assign when_SuperResolutionPart2_l420 = (inpThreshold <= CICC1851_when_SuperResolutionPart2_l419);
  assign when_SuperResolutionPart2_l421 = (inpThreshold <= CICC1851_when_SuperResolutionPart2_l419);
  assign when_SuperResolutionPart2_l422 = (inpThreshold <= CICC1851_when_SuperResolutionPart2_l419);
  assign when_SuperResolutionPart2_l428 = ((inpThreshold <= CICC1851_when_SuperResolutionPart2_l419) && (inpThreshold <= CICC1851_when_SuperResolutionPart2_l428));
  assign when_SuperResolutionPart2_l429 = ((inpThreshold <= CICC1851_when_SuperResolutionPart2_l419) && (inpThreshold <= CICC1851_when_SuperResolutionPart2_l428));
  assign when_SuperResolutionPart2_l430 = (inpThreshold <= CICC1851_when_SuperResolutionPart2_l419);
  assign when_SuperResolutionPart2_l431 = (inpThreshold <= CICC1851_when_SuperResolutionPart2_l419);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_valid = diffStage_controlPipe_fork_io_outputs_0_valid;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_payload_frameStart = diffStage_controlPipe_payload_frameStart;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_payload_rowEnd = diffStage_controlPipe_payload_rowEnd;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_payload_passMode = diffStage_controlPipe_payload_passMode;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_payload_passValid = diffStage_controlPipe_payload_passValid;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceMode = CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceMode;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceValid = CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceValid;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_payload_mainCompare = diffStage_controlPipe_payload_mainCompare;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_payload_counterCompare = diffStage_controlPipe_payload_counterCompare;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_payload_mainDiff = CICC1851_when_SuperResolutionPart2_l419;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_payload_counterDiff = CICC1851_when_SuperResolutionPart2_l428;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceCompValid = CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceCompValid;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceMode = CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceMode;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag = CICC1851_diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_payload_oddValid = diffStage_controlPipe_payload_oddValid;
  assign diffStage_controlPipe_fork_io_outputs_0_translated_ready = (! diffStage_controlPipe_fork_io_outputs_0_translated_rValid);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_valid = (diffStage_controlPipe_fork_io_outputs_0_translated_valid || diffStage_controlPipe_fork_io_outputs_0_translated_rValid);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_frameStart = (diffStage_controlPipe_fork_io_outputs_0_translated_rValid ? diffStage_controlPipe_fork_io_outputs_0_translated_rData_frameStart : diffStage_controlPipe_fork_io_outputs_0_translated_payload_frameStart);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_rowEnd = (diffStage_controlPipe_fork_io_outputs_0_translated_rValid ? diffStage_controlPipe_fork_io_outputs_0_translated_rData_rowEnd : diffStage_controlPipe_fork_io_outputs_0_translated_payload_rowEnd);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_passMode = (diffStage_controlPipe_fork_io_outputs_0_translated_rValid ? diffStage_controlPipe_fork_io_outputs_0_translated_rData_passMode : diffStage_controlPipe_fork_io_outputs_0_translated_payload_passMode);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_passValid = (diffStage_controlPipe_fork_io_outputs_0_translated_rValid ? diffStage_controlPipe_fork_io_outputs_0_translated_rData_passValid : diffStage_controlPipe_fork_io_outputs_0_translated_payload_passValid);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_onceMode = (diffStage_controlPipe_fork_io_outputs_0_translated_rValid ? diffStage_controlPipe_fork_io_outputs_0_translated_rData_onceMode : diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceMode);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_onceValid = (diffStage_controlPipe_fork_io_outputs_0_translated_rValid ? diffStage_controlPipe_fork_io_outputs_0_translated_rData_onceValid : diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceValid);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_mainCompare = (diffStage_controlPipe_fork_io_outputs_0_translated_rValid ? diffStage_controlPipe_fork_io_outputs_0_translated_rData_mainCompare : diffStage_controlPipe_fork_io_outputs_0_translated_payload_mainCompare);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_counterCompare = (diffStage_controlPipe_fork_io_outputs_0_translated_rValid ? diffStage_controlPipe_fork_io_outputs_0_translated_rData_counterCompare : diffStage_controlPipe_fork_io_outputs_0_translated_payload_counterCompare);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_mainDiff = (diffStage_controlPipe_fork_io_outputs_0_translated_rValid ? diffStage_controlPipe_fork_io_outputs_0_translated_rData_mainDiff : diffStage_controlPipe_fork_io_outputs_0_translated_payload_mainDiff);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_counterDiff = (diffStage_controlPipe_fork_io_outputs_0_translated_rValid ? diffStage_controlPipe_fork_io_outputs_0_translated_rData_counterDiff : diffStage_controlPipe_fork_io_outputs_0_translated_payload_counterDiff);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_twiceCompValid = (diffStage_controlPipe_fork_io_outputs_0_translated_rValid ? diffStage_controlPipe_fork_io_outputs_0_translated_rData_twiceCompValid : diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceCompValid);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_twiceMode = (diffStage_controlPipe_fork_io_outputs_0_translated_rValid ? diffStage_controlPipe_fork_io_outputs_0_translated_rData_twiceMode : diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceMode);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_inpValidFlag = (diffStage_controlPipe_fork_io_outputs_0_translated_rValid ? diffStage_controlPipe_fork_io_outputs_0_translated_rData_inpValidFlag : diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag);
  assign diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_oddValid = (diffStage_controlPipe_fork_io_outputs_0_translated_rValid ? diffStage_controlPipe_fork_io_outputs_0_translated_rData_oddValid : diffStage_controlPipe_fork_io_outputs_0_translated_payload_oddValid);
  always @(*) begin
    diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_ready = resultStage_controlPipe_ready;
    if(when_Stream_l368_31) begin
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_31 = (! resultStage_controlPipe_valid);
  assign resultStage_controlPipe_valid = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rValid;
  assign resultStage_controlPipe_payload_frameStart = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_frameStart;
  assign resultStage_controlPipe_payload_rowEnd = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_rowEnd;
  assign resultStage_controlPipe_payload_passMode = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_passMode;
  assign resultStage_controlPipe_payload_passValid = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_passValid;
  assign resultStage_controlPipe_payload_onceMode = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_onceMode;
  assign resultStage_controlPipe_payload_onceValid = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_onceValid;
  assign resultStage_controlPipe_payload_mainCompare = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_mainCompare;
  assign resultStage_controlPipe_payload_counterCompare = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_counterCompare;
  assign resultStage_controlPipe_payload_mainDiff = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_mainDiff;
  assign resultStage_controlPipe_payload_counterDiff = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_counterDiff;
  assign resultStage_controlPipe_payload_twiceCompValid = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_twiceCompValid;
  assign resultStage_controlPipe_payload_twiceMode = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_twiceMode;
  assign resultStage_controlPipe_payload_inpValidFlag = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_inpValidFlag;
  assign resultStage_controlPipe_payload_oddValid = diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_oddValid;
  assign resultStage_pixelStream_valid = diffStage_controlPipe_fork_io_outputs_1_valid;
  always @(*) begin
    resultStage_pixelStream_payload = 8'h0;
    if(diffStage_controlPipe_fork_io_outputs_1_payload_passValid) begin
      if(diffStage_controlPipe_fork_io_outputs_1_payload_passMode) begin
        resultStage_pixelStream_payload = diffStage_mainTwoPixelStream_payload;
      end else begin
        resultStage_pixelStream_payload = diffStage_mainOnePixelStream_payload;
      end
    end
    if(diffStage_controlPipe_fork_io_outputs_1_payload_oddValid) begin
      resultStage_pixelStream_payload = diffStage_oddRowPixelStream_payload;
    end
    if(diffStage_controlPipe_fork_io_outputs_1_payload_onceValid) begin
      case(diffStage_controlPipe_fork_io_outputs_1_payload_onceMode)
        3'b000 : begin
          if(when_SuperResolutionPart2_l451) begin
            resultStage_pixelStream_payload = 8'h0;
          end else begin
            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload[7:0];
          end
        end
        3'b001 : begin
          if(when_SuperResolutionPart2_l455) begin
            resultStage_pixelStream_payload = 8'h0;
          end else begin
            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_2[7:0];
          end
        end
        3'b010 : begin
          if(when_SuperResolutionPart2_l459) begin
            resultStage_pixelStream_payload = 8'h0;
          end else begin
            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_4[7:0];
          end
        end
        3'b011 : begin
          if(when_SuperResolutionPart2_l463) begin
            resultStage_pixelStream_payload = 8'h0;
          end else begin
            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_6[7:0];
          end
        end
        3'b100 : begin
          resultStage_pixelStream_payload = diffStage_mainOnePixelStream_payload;
        end
        3'b101 : begin
          resultStage_pixelStream_payload = diffStage_mainTwoPixelStream_payload;
        end
        default : begin
        end
      endcase
    end
    if(diffStage_controlPipe_fork_io_outputs_1_payload_twiceCompValid) begin
      case(diffStage_controlPipe_fork_io_outputs_1_payload_twiceMode)
        3'b000 : begin
          if(when_SuperResolutionPart2_l474) begin
            resultStage_pixelStream_payload = 8'h0;
          end else begin
            if(when_SuperResolutionPart2_l477) begin
              resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_8[7:0];
            end else begin
              resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_10[7:0];
            end
          end
        end
        3'b001 : begin
          if(when_SuperResolutionPart2_l482) begin
            resultStage_pixelStream_payload = 8'h0;
          end else begin
            if(when_SuperResolutionPart2_l485) begin
              resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_12[7:0];
            end else begin
              resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_14[7:0];
            end
          end
        end
        3'b010 : begin
          resultStage_pixelStream_payload = diffStage_mainTwoPixelStream_payload;
        end
        3'b011 : begin
          if(when_SuperResolutionPart2_l491) begin
            resultStage_pixelStream_payload = 8'h0;
          end else begin
            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_16[7:0];
          end
        end
        3'b100 : begin
          resultStage_pixelStream_payload = diffStage_mainOnePixelStream_payload;
        end
        3'b101 : begin
          if(when_SuperResolutionPart2_l496) begin
            resultStage_pixelStream_payload = 8'h0;
          end else begin
            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_18[7:0];
          end
        end
        default : begin
        end
      endcase
    end
  end

  assign when_SuperResolutionPart2_l451 = (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart2_l455 = (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart2_l459 = (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart2_l463 = (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart2_l474 = ((inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff) && (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff));
  assign when_SuperResolutionPart2_l477 = (diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart2_l482 = ((inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff) && (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff));
  assign when_SuperResolutionPart2_l485 = (diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart2_l491 = (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart2_l496 = (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign resultStage_pixelStream_ready = (! resultStage_pixelStream_rValid);
  assign resultStage_pixelStream_s2mPipe_valid = (resultStage_pixelStream_valid || resultStage_pixelStream_rValid);
  assign resultStage_pixelStream_s2mPipe_payload = (resultStage_pixelStream_rValid ? resultStage_pixelStream_rData : resultStage_pixelStream_payload);
  always @(*) begin
    resultStage_pixelStream_s2mPipe_ready = resultStage_resultStream_ready;
    if(when_Stream_l368_32) begin
      resultStage_pixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_32 = (! resultStage_resultStream_valid);
  assign resultStage_resultStream_valid = resultStage_pixelStream_s2mPipe_rValid;
  assign resultStage_resultStream_payload = resultStage_pixelStream_s2mPipe_rData;
  assign CICC1851_resultStage_mainOnePixelStream_ready_2 = (CICC1851_resultStage_mainOnePixelStream_ready && CICC1851_resultStage_mainOnePixelStream_ready_1);
  assign CICC1851_resultStage_mainOnePixelStream_ready = ((((((resultStage_resultStream_valid && resultStage_mainOnePixelStream_valid) && resultStage_counterOnePixelStream_valid) && resultStage_mainTwoPixelStream_valid) && resultStage_counterTwoPixelStream_valid) && resultStage_controlPipe_valid) && resultStage_oddRowPixelStream_valid);
  assign resultStage_resultStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_mainOnePixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_counterOnePixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_mainTwoPixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_counterTwoPixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_controlPipe_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_oddRowPixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign when_Stream_l438 = ((((! resultStage_controlPipe_payload_passValid) && (! resultStage_controlPipe_payload_onceValid)) && (! resultStage_controlPipe_payload_twiceCompValid)) && (! resultStage_controlPipe_payload_oddValid));
  always @(*) begin
    resultsJoin_valid = CICC1851_resultStage_mainOnePixelStream_ready;
    if(when_Stream_l438) begin
      resultsJoin_valid = 1'b0;
    end
  end

  always @(*) begin
    CICC1851_resultStage_mainOnePixelStream_ready_1 = resultsJoin_ready;
    if(when_Stream_l438) begin
      CICC1851_resultStage_mainOnePixelStream_ready_1 = 1'b1;
    end
  end

  assign pixelsStream_valid = resultsJoin_valid;
  assign resultsJoin_ready = pixelsStream_ready;
  assign pixelsStream_payload_pixel = resultStage_resultStream_payload;
  assign pixelsStream_payload_frameStart = resultStage_controlPipe_payload_frameStart;
  assign pixelsStream_payload_rowEnd = resultStage_controlPipe_payload_rowEnd;
  assign pixelsStream_payload_inpValid = resultStage_controlPipe_payload_inpValidFlag;
  assign pixelsStream_ready = (! pixelsStream_rValid);
  assign pixelsStream_s2mPipe_valid = (pixelsStream_valid || pixelsStream_rValid);
  assign pixelsStream_s2mPipe_payload_pixel = (pixelsStream_rValid ? pixelsStream_rData_pixel : pixelsStream_payload_pixel);
  assign pixelsStream_s2mPipe_payload_frameStart = (pixelsStream_rValid ? pixelsStream_rData_frameStart : pixelsStream_payload_frameStart);
  assign pixelsStream_s2mPipe_payload_rowEnd = (pixelsStream_rValid ? pixelsStream_rData_rowEnd : pixelsStream_payload_rowEnd);
  assign pixelsStream_s2mPipe_payload_inpValid = (pixelsStream_rValid ? pixelsStream_rData_inpValid : pixelsStream_payload_inpValid);
  always @(*) begin
    pixelsStream_s2mPipe_ready = pixelsStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_33) begin
      pixelsStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_33 = (! pixelsStream_s2mPipe_m2sPipe_valid);
  assign pixelsStream_s2mPipe_m2sPipe_valid = pixelsStream_s2mPipe_rValid;
  assign pixelsStream_s2mPipe_m2sPipe_payload_pixel = pixelsStream_s2mPipe_rData_pixel;
  assign pixelsStream_s2mPipe_m2sPipe_payload_frameStart = pixelsStream_s2mPipe_rData_frameStart;
  assign pixelsStream_s2mPipe_m2sPipe_payload_rowEnd = pixelsStream_s2mPipe_rData_rowEnd;
  assign pixelsStream_s2mPipe_m2sPipe_payload_inpValid = pixelsStream_s2mPipe_rData_inpValid;
  assign pixelsStream_s2mPipe_m2sPipe_ready = pixelsOut_ready;
  assign controlStateMachine_wantExit = 1'b0;
  always @(*) begin
    controlStateMachine_wantStart = 1'b0;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_1_HOLD : begin
      end
      controlStateMachine_enumDef_1_PASS : begin
      end
      controlStateMachine_enumDef_1_ONCE : begin
      end
      controlStateMachine_enumDef_1_TWICE : begin
      end
      default : begin
        controlStateMachine_wantStart = 1'b1;
      end
    endcase
  end

  assign controlStateMachine_wantKill = 1'b0;
  assign when_SuperResolutionPart2_l761 = (((currentState == 3'b010) || (currentState == 3'b011)) || (currentState == 3'b100));
  assign controlStream_fire_4 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart2_l763 = (controlStream_fire_4 && (CICC1851_when_SuperResolutionPart2_l763 == CICC1851_when_SuperResolutionPart2_l763_1));
  assign controlStream_fire_5 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart2_l764 = ((outReachRowEnd && (CICC1851_when_SuperResolutionPart2_l764 == CICC1851_when_SuperResolutionPart2_l764_1)) && controlStream_fire_5);
  assign controlStream_fire_6 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart2_l766 = (controlStream_fire_6 && outReachRowEnd);
  assign controlStream_fire_7 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart2_l783 = (CICC1851_when_SuperResolutionPart2_l783 == 12'h0);
  assign when_SuperResolutionPart2_l785 = (CICC1851_when_SuperResolutionPart2_l785 == 12'h001);
  assign when_SuperResolutionPart2_l787 = (CICC1851_when_SuperResolutionPart2_l787 == 12'h002);
  assign when_SuperResolutionPart2_l789 = (CICC1851_when_SuperResolutionPart2_l789 == 12'h003);
  assign when_SuperResolutionPart2_l793 = (CICC1851_when_SuperResolutionPart2_l793 == 12'h0);
  assign when_SuperResolutionPart2_l796 = (CICC1851_when_SuperResolutionPart2_l796 == 12'h001);
  assign when_SuperResolutionPart2_l799 = (CICC1851_when_SuperResolutionPart2_l799 == 12'h002);
  assign when_SuperResolutionPart2_l802 = (CICC1851_when_SuperResolutionPart2_l802 == 12'h003);
  always @(*) begin
    controlStateMachine_stateNext = controlStateMachine_stateReg;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_1_HOLD : begin
        if(zeroInFourOutRow) begin
          if(passPixels_fire_13) begin
            if(threeInFourOutPixelAddr) begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_1_ONCE;
            end else begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_1_PASS;
            end
          end
        end else begin
          if(twoInFourOutRow) begin
            if(passPixels_fire_14) begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_1_PASS;
            end
          end else begin
            if(threeInFourOutRow) begin
              if(passPixels_fire_15) begin
                if(threeInFourOutPixelAddr) begin
                  if(willHoldToTwice) begin
                    controlStateMachine_stateNext = controlStateMachine_enumDef_1_TWICE;
                  end
                end else begin
                  controlStateMachine_stateNext = controlStateMachine_enumDef_1_ONCE;
                end
              end
            end
          end
        end
      end
      controlStateMachine_enumDef_1_PASS : begin
        if(controlStream_fire_8) begin
          if(oneInFourOutPixelAddr) begin
            if(oneInFourOutRow) begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_1_PASS;
            end else begin
              if(twoInFourOutRow) begin
                if(when_SuperResolutionPart2_l573) begin
                  controlStateMachine_stateNext = controlStateMachine_enumDef_1_HOLD;
                end else begin
                  controlStateMachine_stateNext = controlStateMachine_enumDef_1_PASS;
                end
              end else begin
                if(when_SuperResolutionPart2_l578) begin
                  controlStateMachine_stateNext = controlStateMachine_enumDef_1_HOLD;
                end else begin
                  controlStateMachine_stateNext = controlStateMachine_enumDef_1_PASS;
                end
              end
            end
          end else begin
            if(twoInFourOutPixelAddr) begin
              if(oneInFourOutRow) begin
                controlStateMachine_stateNext = controlStateMachine_enumDef_1_ONCE;
              end else begin
                if(twoInFourOutRow) begin
                  controlStateMachine_stateNext = controlStateMachine_enumDef_1_ONCE;
                end else begin
                  if(when_SuperResolutionPart2_l590) begin
                    controlStateMachine_stateNext = controlStateMachine_enumDef_1_HOLD;
                  end else begin
                    controlStateMachine_stateNext = controlStateMachine_enumDef_1_ONCE;
                  end
                end
              end
            end else begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_1_PASS;
            end
          end
        end
      end
      controlStateMachine_enumDef_1_ONCE : begin
        if(controlStream_fire_10) begin
          if(zeroInFourOutRow) begin
            controlStateMachine_stateNext = controlStateMachine_enumDef_1_PASS;
          end else begin
            if(oneInFourOutRow) begin
              if(when_SuperResolutionPart2_l642) begin
                controlStateMachine_stateNext = controlStateMachine_enumDef_1_HOLD;
              end else begin
                controlStateMachine_stateNext = controlStateMachine_enumDef_1_PASS;
              end
            end else begin
              if(twoInFourOutRow) begin
                if(outReachRowEnd) begin
                  if(when_SuperResolutionPart2_l647) begin
                    controlStateMachine_stateNext = controlStateMachine_enumDef_1_HOLD;
                  end else begin
                    controlStateMachine_stateNext = controlStateMachine_enumDef_1_ONCE;
                  end
                end else begin
                  controlStateMachine_stateNext = controlStateMachine_enumDef_1_PASS;
                end
              end else begin
                if(twoInFourOutPixelAddr) begin
                  if(when_SuperResolutionPart2_l653) begin
                    controlStateMachine_stateNext = controlStateMachine_enumDef_1_HOLD;
                  end else begin
                    controlStateMachine_stateNext = controlStateMachine_enumDef_1_TWICE;
                  end
                end else begin
                  controlStateMachine_stateNext = controlStateMachine_enumDef_1_ONCE;
                end
              end
            end
          end
        end
      end
      controlStateMachine_enumDef_1_TWICE : begin
        if(controlStream_fire_11) begin
          if(outReachRowEnd) begin
            if(outReachFinalRow) begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_1_HOLD;
            end else begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_1_PASS;
            end
          end else begin
            controlStateMachine_stateNext = controlStateMachine_enumDef_1_ONCE;
          end
        end
      end
      default : begin
      end
    endcase
    if(controlStateMachine_wantStart) begin
      controlStateMachine_stateNext = controlStateMachine_enumDef_1_HOLD;
    end
    if(controlStateMachine_wantKill) begin
      controlStateMachine_stateNext = controlStateMachine_enumDef_1_BOOT;
    end
  end

  assign passPixels_fire_13 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_14 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_15 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_16 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart2_l560 = (CICC1851_when_SuperResolutionPart2_l560 == CICC1851_when_SuperResolutionPart2_l560_1);
  assign controlStream_fire_8 = (controlStream_valid && controlStream_ready);
  assign passPixels_fire_17 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart2_l573 = ((((oddBufferRow && (! holdBuffer)) && willPassToHoldCaseOne) && (! passPixels_fire_17)) && (! bufferReuse));
  assign passPixels_fire_18 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart2_l578 = (((((! oddBufferRow) && (! holdBuffer)) && willPassToHoldCaseOne) && (! passPixels_fire_18)) && (! bufferReuse));
  assign when_SuperResolutionPart2_l585 = ((oddBufferRow && (! holdBuffer)) && (! bufferReachRowEnd));
  assign when_SuperResolutionPart2_l588 = (((! oddBufferRow) && (! bufferReuse)) && (! bufferReachRowEnd));
  assign passPixels_fire_19 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart2_l590 = (((((! oddBufferRow) && (! holdBuffer)) && (! bufferReuse)) && (willPassToHoldCaseTwo || holdWillPassToHoldCaseTwo)) && (! passPixels_fire_19));
  assign when_SuperResolutionPart2_l602 = (poping && (CICC1851_when_SuperResolutionPart2_l602 == CICC1851_when_SuperResolutionPart2_l602_1));
  assign when_SuperResolutionPart2_l603 = (pushAndPoping && (CICC1851_when_SuperResolutionPart2_l603 == CICC1851_when_SuperResolutionPart2_l603_1));
  assign when_SuperResolutionPart2_l605 = (poping && (CICC1851_when_SuperResolutionPart2_l605 == CICC1851_when_SuperResolutionPart2_l605_1));
  assign when_SuperResolutionPart2_l606 = (pushAndPoping && (CICC1851_when_SuperResolutionPart2_l606 == CICC1851_when_SuperResolutionPart2_l606_1));
  assign when_SuperResolutionPart2_l609 = (CICC1851_when_SuperResolutionPart2_l609 == 12'h0);
  assign controlStream_fire_9 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart2_l630 = (frameStart && controlStream_fire_9);
  assign controlStream_fire_10 = (controlStream_valid && controlStream_ready);
  assign passPixels_fire_20 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart2_l642 = (((outReachRowEnd && willOnceToHoldCaseOne) && (bufferWAddr_value == 11'h0)) && (! passPixels_fire_20));
  assign passPixels_fire_21 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart2_l647 = (((bufferWAddr_value == 11'h0) && (! passPixels_fire_21)) && willOnceToHoldCaseTwo);
  assign passPixels_fire_22 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart2_l653 = ((((! oddBufferRow) && willOnceToHoldCaseThree) && (! passPixels_fire_22)) && (! bufferReuse));
  assign passPixels_fire_23 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart2_l662 = (passPixels_fire_23 && bufferReachRowEnd);
  assign when_SuperResolutionPart2_l667 = (poping && (CICC1851_when_SuperResolutionPart2_l667 == CICC1851_when_SuperResolutionPart2_l667_2));
  assign when_SuperResolutionPart2_l668 = (pushAndPoping && (CICC1851_when_SuperResolutionPart2_l668 == CICC1851_when_SuperResolutionPart2_l668_1));
  assign controlStream_fire_11 = (controlStream_valid && controlStream_ready);
  assign currentState = controlStateMachine_stateReg;
  always @(posedge clk or negedge resetn) begin
    if(!resetn) begin
      inpTwoDone <= 1'b0;
      readDone <= 1'b0;
      startRead <= 1'b0;
      slaveStart <= 1'b0;
      frameStart <= 1'b0;
      inpThreshold <= 8'h80;
      bmpWidth <= 10'h3c0;
      bmpHeight <= 10'h21c;
      holdBuffer <= 1'b0;
      writeDone <= 1'b0;
      bufferRowCount_value <= 11'h0;
      bufferReuse <= 1'b0;
      bufferEnable <= 1'b0;
      bufferSwitch <= 2'b00;
      nextRowBuffer <= 1'b1;
      bufferWAddr_value <= 11'h0;
      outPixelAddr_value <= 12'h0;
      outRowCount_value <= 12'h0;
      alreadySendRow_value <= 12'h0;
      alreadySendCountInRow_value <= 12'h0;
      alreadyReachRowEnd <= 1'b0;
      alreadyReachFinalRow <= 1'b0;
      outReachRowEnd <= 1'b0;
      outReachFinalRow <= 1'b0;
      bufferReachRowEnd <= 1'b0;
      bufferReachFinalRow <= 1'b0;
      oddBufferRow <= 1'b0;
      zeroInFourOutPixelAddr <= 1'b1;
      oneInFourOutPixelAddr <= 1'b0;
      twoInFourOutPixelAddr <= 1'b0;
      threeInFourOutPixelAddr <= 1'b0;
      zeroInFourOutRow <= 1'b1;
      oneInFourOutRow <= 1'b0;
      twoInFourOutRow <= 1'b0;
      threeInFourOutRow <= 1'b0;
      willHoldToTwice <= 1'b0;
      willPassToHoldCaseOne <= 1'b0;
      willPassToHoldCaseTwo <= 1'b0;
      holdWillPassToHoldCaseTwo <= 1'b0;
      willOnceToHoldCaseOne <= 1'b0;
      willOnceToHoldCaseTwo <= 1'b0;
      willOnceToHoldCaseThree <= 1'b0;
      pixelsIn_rValid <= 1'b0;
      pixelsIn_s2mPipe_rValid <= 1'b0;
      mainAddrOneStream_rValid <= 1'b0;
      mainAddrOneStream_s2mPipe_rValid <= 1'b0;
      CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_mainOnePixelStream_valid <= 1'b0;
      counterAddrOneStream_rValid <= 1'b0;
      counterAddrOneStream_s2mPipe_rValid <= 1'b0;
      CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_counterOnePixelStream_valid <= 1'b0;
      mainAddrTwoStream_rValid <= 1'b0;
      mainAddrTwoStream_s2mPipe_rValid <= 1'b0;
      CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_mainTwoPixelStream_valid <= 1'b0;
      counterAddrTwoStream_rValid <= 1'b0;
      counterAddrTwoStream_s2mPipe_rValid <= 1'b0;
      CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_counterTwoPixelStream_valid <= 1'b0;
      oddAddrStream_rValid <= 1'b0;
      oddAddrStream_s2mPipe_rValid <= 1'b0;
      CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_oddRowPixelStream_valid <= 1'b0;
      controlStream_rValid <= 1'b0;
      controlStream_s2mPipe_rValid <= 1'b0;
      controlStream_s2mPipe_m2sPipe_rValid <= 1'b0;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rValid <= 1'b0;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rValid <= 1'b0;
      readStage_mainOnePixelStream_rValid <= 1'b0;
      readStage_mainOnePixelStream_s2mPipe_rValid <= 1'b0;
      readStage_counterOnePixelStream_rValid <= 1'b0;
      readStage_counterOnePixelStream_s2mPipe_rValid <= 1'b0;
      readStage_mainTwoPixelStream_rValid <= 1'b0;
      readStage_mainTwoPixelStream_s2mPipe_rValid <= 1'b0;
      readStage_counterTwoPixelStream_rValid <= 1'b0;
      readStage_counterTwoPixelStream_s2mPipe_rValid <= 1'b0;
      readStage_oddRowPixelStream_rValid <= 1'b0;
      readStage_oddRowPixelStream_s2mPipe_rValid <= 1'b0;
      readStage_controlPipe_translated_rValid <= 1'b0;
      readStage_controlPipe_translated_s2mPipe_rValid <= 1'b0;
      compareStage_mainOnePixelStream_rValid <= 1'b0;
      compareStage_mainOnePixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_counterOnePixelStream_rValid <= 1'b0;
      compareStage_counterOnePixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_mainTwoPixelStream_rValid <= 1'b0;
      compareStage_mainTwoPixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_counterTwoPixelStream_rValid <= 1'b0;
      compareStage_counterTwoPixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_oddRowPixelStream_rValid <= 1'b0;
      compareStage_oddRowPixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_controlPipe_translated_rValid <= 1'b0;
      compareStage_controlPipe_translated_s2mPipe_rValid <= 1'b0;
      diffStage_mainOnePixelStream_rValid <= 1'b0;
      diffStage_mainOnePixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_counterOnePixelStream_rValid <= 1'b0;
      diffStage_counterOnePixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_mainTwoPixelStream_rValid <= 1'b0;
      diffStage_mainTwoPixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_counterTwoPixelStream_rValid <= 1'b0;
      diffStage_counterTwoPixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_oddRowPixelStream_rValid <= 1'b0;
      diffStage_oddRowPixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_controlPipe_fork_io_outputs_0_translated_rValid <= 1'b0;
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rValid <= 1'b0;
      resultStage_pixelStream_rValid <= 1'b0;
      resultStage_pixelStream_s2mPipe_rValid <= 1'b0;
      pixelsStream_rValid <= 1'b0;
      pixelsStream_s2mPipe_rValid <= 1'b0;
      controlStateMachine_stateReg <= controlStateMachine_enumDef_1_BOOT;
    end else begin
      if(when_SuperResolutionPart2_l40) begin
        inpTwoDone <= 1'b0;
      end
      if(when_SuperResolutionPart2_l43) begin
        readDone <= 1'b0;
      end
      if(when_SuperResolutionPart2_l46) begin
        startRead <= 1'b1;
      end
      if(when_SuperResolutionPart2_l46_1) begin
        startRead <= 1'b0;
      end
      if(when_SuperResolutionPart2_l49) begin
        slaveStart <= 1'b1;
      end
      if(when_SuperResolutionPart2_l49_1) begin
        slaveStart <= 1'b0;
      end
      inpThreshold <= thresholdIn;
      bmpWidth <= widthIn;
      bmpHeight <= heightIn;
      if(when_SuperResolutionPart2_l64) begin
        holdBuffer <= 1'b0;
      end
      if(when_SuperResolutionPart2_l67) begin
        writeDone <= 1'b0;
      end
      bufferRowCount_value <= bufferRowCount_valueNext;
      if(inpTwoDone) begin
        bufferReuse <= 1'b0;
      end
      if(when_SuperResolutionPart2_l76) begin
        bufferEnable <= 1'b1;
      end
      if(when_SuperResolutionPart2_l76_1) begin
        bufferEnable <= 1'b0;
      end
      if(when_SuperResolutionPart2_l82) begin
        nextRowBuffer <= 1'b1;
      end
      bufferWAddr_value <= bufferWAddr_valueNext;
      outPixelAddr_value <= outPixelAddr_valueNext;
      outRowCount_value <= outRowCount_valueNext;
      alreadySendRow_value <= alreadySendRow_valueNext;
      alreadySendCountInRow_value <= alreadySendCountInRow_valueNext;
      if(when_SuperResolutionPart2_l106) begin
        oddBufferRow <= 1'b0;
      end
      if(when_SuperResolutionPart2_l108) begin
        zeroInFourOutPixelAddr <= 1'b1;
      end
      if(when_SuperResolutionPart2_l109) begin
        oneInFourOutPixelAddr <= 1'b0;
      end
      if(when_SuperResolutionPart2_l110) begin
        twoInFourOutPixelAddr <= 1'b0;
      end
      if(when_SuperResolutionPart2_l111) begin
        threeInFourOutPixelAddr <= 1'b0;
      end
      if(when_SuperResolutionPart2_l113) begin
        zeroInFourOutRow <= 1'b1;
      end
      if(when_SuperResolutionPart2_l114) begin
        oneInFourOutRow <= 1'b0;
      end
      if(when_SuperResolutionPart2_l115) begin
        twoInFourOutRow <= 1'b0;
      end
      if(when_SuperResolutionPart2_l116) begin
        threeInFourOutRow <= 1'b0;
      end
      if(when_SuperResolutionPart2_l120) begin
        willHoldToTwice <= 1'b0;
      end
      if(when_SuperResolutionPart2_l121) begin
        willPassToHoldCaseOne <= 1'b0;
      end
      if(when_SuperResolutionPart2_l122) begin
        willPassToHoldCaseTwo <= 1'b0;
      end
      if(when_SuperResolutionPart2_l123) begin
        holdWillPassToHoldCaseTwo <= 1'b0;
      end
      if(when_SuperResolutionPart2_l124) begin
        willOnceToHoldCaseOne <= 1'b0;
      end
      if(when_SuperResolutionPart2_l125) begin
        willOnceToHoldCaseTwo <= 1'b0;
      end
      if(when_SuperResolutionPart2_l126) begin
        willOnceToHoldCaseThree <= 1'b0;
      end
      if(when_SuperResolutionPart2_l134) begin
        bufferSwitch <= 2'b00;
      end
      if(pixelsIn_valid) begin
        pixelsIn_rValid <= 1'b1;
      end
      if(pixelsIn_s2mPipe_ready) begin
        pixelsIn_rValid <= 1'b0;
      end
      if(pixelsIn_s2mPipe_ready) begin
        pixelsIn_s2mPipe_rValid <= pixelsIn_s2mPipe_valid;
      end
      if(when_SuperResolutionPart2_l181) begin
        bufferReachRowEnd <= 1'b1;
      end
      if(when_SuperResolutionPart2_l182) begin
        bufferReachFinalRow <= 1'b1;
      end
      if(when_SuperResolutionPart2_l185) begin
        if(bufferReachFinalRow) begin
          bufferReachRowEnd <= 1'b0;
          bufferReachFinalRow <= 1'b0;
          bufferReuse <= 1'b1;
        end else begin
          bufferReachRowEnd <= 1'b0;
        end
        if(when_SuperResolutionPart2_l195) begin
          oddBufferRow <= 1'b1;
        end else begin
          oddBufferRow <= 1'b0;
        end
      end
      if(when_SuperResolutionPart2_l200) begin
        if(when_SuperResolutionPart2_l201) begin
          bufferSwitch <= 2'b01;
        end else begin
          if(nextRowBuffer) begin
            bufferSwitch <= (bufferSwitch + 2'b01);
          end else begin
            bufferSwitch <= (bufferSwitch - 2'b01);
          end
        end
      end
      if(when_SuperResolutionPart2_l207) begin
        if(when_SuperResolutionPart2_l208) begin
          holdBuffer <= 1'b1;
          bufferEnable <= 1'b0;
        end
        if(when_SuperResolutionPart2_l212) begin
          writeDone <= 1'b1;
          bufferEnable <= 1'b0;
        end
      end
      if(when_SuperResolutionPart2_l218) begin
        holdBuffer <= 1'b0;
        if(when_SuperResolutionPart2_l220) begin
          nextRowBuffer <= (! nextRowBuffer);
        end
      end
      if(when_SuperResolutionPart2_l224) begin
        frameStart <= 1'b1;
      end
      if(when_SuperResolutionPart2_l234) begin
        alreadyReachRowEnd <= 1'b1;
      end
      if(when_SuperResolutionPart2_l235) begin
        alreadyReachFinalRow <= 1'b1;
      end
      if(pixelsOut_fire_2) begin
        if(alreadyReachRowEnd) begin
          alreadyReachRowEnd <= 1'b0;
          if(alreadyReachFinalRow) begin
            alreadyReachFinalRow <= 1'b0;
          end
        end
      end
      if(when_SuperResolutionPart2_l246) begin
        inpTwoDone <= 1'b1;
      end
      if(mainAddrOneStream_valid) begin
        mainAddrOneStream_rValid <= 1'b1;
      end
      if(mainAddrOneStream_s2mPipe_ready) begin
        mainAddrOneStream_rValid <= 1'b0;
      end
      if(mainAddrOneStream_s2mPipe_ready) begin
        mainAddrOneStream_s2mPipe_rValid <= mainAddrOneStream_s2mPipe_valid;
      end
      if(CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(mainAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_2 <= mainAddrOneStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_1) begin
        CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_1) begin
        CICC1851_readStage_mainOnePixelStream_valid <= (CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready || CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_3);
      end
      if(counterAddrOneStream_valid) begin
        counterAddrOneStream_rValid <= 1'b1;
      end
      if(counterAddrOneStream_s2mPipe_ready) begin
        counterAddrOneStream_rValid <= 1'b0;
      end
      if(counterAddrOneStream_s2mPipe_ready) begin
        counterAddrOneStream_s2mPipe_rValid <= counterAddrOneStream_s2mPipe_valid;
      end
      if(CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(counterAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_2 <= counterAddrOneStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_2) begin
        CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_2) begin
        CICC1851_readStage_counterOnePixelStream_valid <= (CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready || CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_3);
      end
      if(mainAddrTwoStream_valid) begin
        mainAddrTwoStream_rValid <= 1'b1;
      end
      if(mainAddrTwoStream_s2mPipe_ready) begin
        mainAddrTwoStream_rValid <= 1'b0;
      end
      if(mainAddrTwoStream_s2mPipe_ready) begin
        mainAddrTwoStream_s2mPipe_rValid <= mainAddrTwoStream_s2mPipe_valid;
      end
      if(CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(mainAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= mainAddrTwoStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_3) begin
        CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_3) begin
        CICC1851_readStage_mainTwoPixelStream_valid <= (CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready || CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_3);
      end
      if(counterAddrTwoStream_valid) begin
        counterAddrTwoStream_rValid <= 1'b1;
      end
      if(counterAddrTwoStream_s2mPipe_ready) begin
        counterAddrTwoStream_rValid <= 1'b0;
      end
      if(counterAddrTwoStream_s2mPipe_ready) begin
        counterAddrTwoStream_s2mPipe_rValid <= counterAddrTwoStream_s2mPipe_valid;
      end
      if(CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(counterAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= counterAddrTwoStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_4) begin
        CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_4) begin
        CICC1851_readStage_counterTwoPixelStream_valid <= (CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready || CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_3);
      end
      if(oddAddrStream_valid) begin
        oddAddrStream_rValid <= 1'b1;
      end
      if(oddAddrStream_s2mPipe_ready) begin
        oddAddrStream_rValid <= 1'b0;
      end
      if(oddAddrStream_s2mPipe_ready) begin
        oddAddrStream_s2mPipe_rValid <= oddAddrStream_s2mPipe_valid;
      end
      if(CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(oddAddrStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_2 <= oddAddrStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_5) begin
        CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_5) begin
        CICC1851_readStage_oddRowPixelStream_valid <= (CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready || CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_3);
      end
      if(controlStream_valid) begin
        controlStream_rValid <= 1'b1;
      end
      if(controlStream_s2mPipe_ready) begin
        controlStream_rValid <= 1'b0;
      end
      if(controlStream_s2mPipe_ready) begin
        controlStream_s2mPipe_rValid <= controlStream_s2mPipe_valid;
      end
      if(controlStream_s2mPipe_m2sPipe_ready) begin
        controlStream_s2mPipe_m2sPipe_rValid <= controlStream_s2mPipe_m2sPipe_valid;
      end
      if(controlStream_s2mPipe_m2sPipe_m2sPipe_valid) begin
        controlStream_s2mPipe_m2sPipe_m2sPipe_rValid <= 1'b1;
      end
      if(controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready) begin
        controlStream_s2mPipe_m2sPipe_m2sPipe_rValid <= 1'b0;
      end
      if(controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready) begin
        controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_valid;
      end
      if(readStage_mainOnePixelStream_valid) begin
        readStage_mainOnePixelStream_rValid <= 1'b1;
      end
      if(readStage_mainOnePixelStream_s2mPipe_ready) begin
        readStage_mainOnePixelStream_rValid <= 1'b0;
      end
      if(readStage_mainOnePixelStream_s2mPipe_ready) begin
        readStage_mainOnePixelStream_s2mPipe_rValid <= readStage_mainOnePixelStream_s2mPipe_valid;
      end
      if(readStage_counterOnePixelStream_valid) begin
        readStage_counterOnePixelStream_rValid <= 1'b1;
      end
      if(readStage_counterOnePixelStream_s2mPipe_ready) begin
        readStage_counterOnePixelStream_rValid <= 1'b0;
      end
      if(readStage_counterOnePixelStream_s2mPipe_ready) begin
        readStage_counterOnePixelStream_s2mPipe_rValid <= readStage_counterOnePixelStream_s2mPipe_valid;
      end
      if(readStage_mainTwoPixelStream_valid) begin
        readStage_mainTwoPixelStream_rValid <= 1'b1;
      end
      if(readStage_mainTwoPixelStream_s2mPipe_ready) begin
        readStage_mainTwoPixelStream_rValid <= 1'b0;
      end
      if(readStage_mainTwoPixelStream_s2mPipe_ready) begin
        readStage_mainTwoPixelStream_s2mPipe_rValid <= readStage_mainTwoPixelStream_s2mPipe_valid;
      end
      if(readStage_counterTwoPixelStream_valid) begin
        readStage_counterTwoPixelStream_rValid <= 1'b1;
      end
      if(readStage_counterTwoPixelStream_s2mPipe_ready) begin
        readStage_counterTwoPixelStream_rValid <= 1'b0;
      end
      if(readStage_counterTwoPixelStream_s2mPipe_ready) begin
        readStage_counterTwoPixelStream_s2mPipe_rValid <= readStage_counterTwoPixelStream_s2mPipe_valid;
      end
      if(readStage_oddRowPixelStream_valid) begin
        readStage_oddRowPixelStream_rValid <= 1'b1;
      end
      if(readStage_oddRowPixelStream_s2mPipe_ready) begin
        readStage_oddRowPixelStream_rValid <= 1'b0;
      end
      if(readStage_oddRowPixelStream_s2mPipe_ready) begin
        readStage_oddRowPixelStream_s2mPipe_rValid <= readStage_oddRowPixelStream_s2mPipe_valid;
      end
      if(readStage_controlPipe_translated_valid) begin
        readStage_controlPipe_translated_rValid <= 1'b1;
      end
      if(readStage_controlPipe_translated_s2mPipe_ready) begin
        readStage_controlPipe_translated_rValid <= 1'b0;
      end
      if(readStage_controlPipe_translated_s2mPipe_ready) begin
        readStage_controlPipe_translated_s2mPipe_rValid <= readStage_controlPipe_translated_s2mPipe_valid;
      end
      if(compareStage_mainOnePixelStream_valid) begin
        compareStage_mainOnePixelStream_rValid <= 1'b1;
      end
      if(compareStage_mainOnePixelStream_s2mPipe_ready) begin
        compareStage_mainOnePixelStream_rValid <= 1'b0;
      end
      if(compareStage_mainOnePixelStream_s2mPipe_ready) begin
        compareStage_mainOnePixelStream_s2mPipe_rValid <= compareStage_mainOnePixelStream_s2mPipe_valid;
      end
      if(compareStage_counterOnePixelStream_valid) begin
        compareStage_counterOnePixelStream_rValid <= 1'b1;
      end
      if(compareStage_counterOnePixelStream_s2mPipe_ready) begin
        compareStage_counterOnePixelStream_rValid <= 1'b0;
      end
      if(compareStage_counterOnePixelStream_s2mPipe_ready) begin
        compareStage_counterOnePixelStream_s2mPipe_rValid <= compareStage_counterOnePixelStream_s2mPipe_valid;
      end
      if(compareStage_mainTwoPixelStream_valid) begin
        compareStage_mainTwoPixelStream_rValid <= 1'b1;
      end
      if(compareStage_mainTwoPixelStream_s2mPipe_ready) begin
        compareStage_mainTwoPixelStream_rValid <= 1'b0;
      end
      if(compareStage_mainTwoPixelStream_s2mPipe_ready) begin
        compareStage_mainTwoPixelStream_s2mPipe_rValid <= compareStage_mainTwoPixelStream_s2mPipe_valid;
      end
      if(compareStage_counterTwoPixelStream_valid) begin
        compareStage_counterTwoPixelStream_rValid <= 1'b1;
      end
      if(compareStage_counterTwoPixelStream_s2mPipe_ready) begin
        compareStage_counterTwoPixelStream_rValid <= 1'b0;
      end
      if(compareStage_counterTwoPixelStream_s2mPipe_ready) begin
        compareStage_counterTwoPixelStream_s2mPipe_rValid <= compareStage_counterTwoPixelStream_s2mPipe_valid;
      end
      if(compareStage_oddRowPixelStream_valid) begin
        compareStage_oddRowPixelStream_rValid <= 1'b1;
      end
      if(compareStage_oddRowPixelStream_s2mPipe_ready) begin
        compareStage_oddRowPixelStream_rValid <= 1'b0;
      end
      if(compareStage_oddRowPixelStream_s2mPipe_ready) begin
        compareStage_oddRowPixelStream_s2mPipe_rValid <= compareStage_oddRowPixelStream_s2mPipe_valid;
      end
      if(compareStage_controlPipe_translated_valid) begin
        compareStage_controlPipe_translated_rValid <= 1'b1;
      end
      if(compareStage_controlPipe_translated_s2mPipe_ready) begin
        compareStage_controlPipe_translated_rValid <= 1'b0;
      end
      if(compareStage_controlPipe_translated_s2mPipe_ready) begin
        compareStage_controlPipe_translated_s2mPipe_rValid <= compareStage_controlPipe_translated_s2mPipe_valid;
      end
      if(diffStage_mainOnePixelStream_valid) begin
        diffStage_mainOnePixelStream_rValid <= 1'b1;
      end
      if(diffStage_mainOnePixelStream_s2mPipe_ready) begin
        diffStage_mainOnePixelStream_rValid <= 1'b0;
      end
      if(diffStage_mainOnePixelStream_s2mPipe_ready) begin
        diffStage_mainOnePixelStream_s2mPipe_rValid <= diffStage_mainOnePixelStream_s2mPipe_valid;
      end
      if(diffStage_counterOnePixelStream_valid) begin
        diffStage_counterOnePixelStream_rValid <= 1'b1;
      end
      if(diffStage_counterOnePixelStream_s2mPipe_ready) begin
        diffStage_counterOnePixelStream_rValid <= 1'b0;
      end
      if(diffStage_counterOnePixelStream_s2mPipe_ready) begin
        diffStage_counterOnePixelStream_s2mPipe_rValid <= diffStage_counterOnePixelStream_s2mPipe_valid;
      end
      if(diffStage_mainTwoPixelStream_valid) begin
        diffStage_mainTwoPixelStream_rValid <= 1'b1;
      end
      if(diffStage_mainTwoPixelStream_s2mPipe_ready) begin
        diffStage_mainTwoPixelStream_rValid <= 1'b0;
      end
      if(diffStage_mainTwoPixelStream_s2mPipe_ready) begin
        diffStage_mainTwoPixelStream_s2mPipe_rValid <= diffStage_mainTwoPixelStream_s2mPipe_valid;
      end
      if(diffStage_counterTwoPixelStream_valid) begin
        diffStage_counterTwoPixelStream_rValid <= 1'b1;
      end
      if(diffStage_counterTwoPixelStream_s2mPipe_ready) begin
        diffStage_counterTwoPixelStream_rValid <= 1'b0;
      end
      if(diffStage_counterTwoPixelStream_s2mPipe_ready) begin
        diffStage_counterTwoPixelStream_s2mPipe_rValid <= diffStage_counterTwoPixelStream_s2mPipe_valid;
      end
      if(diffStage_oddRowPixelStream_valid) begin
        diffStage_oddRowPixelStream_rValid <= 1'b1;
      end
      if(diffStage_oddRowPixelStream_s2mPipe_ready) begin
        diffStage_oddRowPixelStream_rValid <= 1'b0;
      end
      if(diffStage_oddRowPixelStream_s2mPipe_ready) begin
        diffStage_oddRowPixelStream_s2mPipe_rValid <= diffStage_oddRowPixelStream_s2mPipe_valid;
      end
      if(diffStage_controlPipe_fork_io_outputs_0_translated_valid) begin
        diffStage_controlPipe_fork_io_outputs_0_translated_rValid <= 1'b1;
      end
      if(diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_ready) begin
        diffStage_controlPipe_fork_io_outputs_0_translated_rValid <= 1'b0;
      end
      if(diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_ready) begin
        diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rValid <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_valid;
      end
      if(resultStage_pixelStream_valid) begin
        resultStage_pixelStream_rValid <= 1'b1;
      end
      if(resultStage_pixelStream_s2mPipe_ready) begin
        resultStage_pixelStream_rValid <= 1'b0;
      end
      if(resultStage_pixelStream_s2mPipe_ready) begin
        resultStage_pixelStream_s2mPipe_rValid <= resultStage_pixelStream_s2mPipe_valid;
      end
      if(pixelsStream_valid) begin
        pixelsStream_rValid <= 1'b1;
      end
      if(pixelsStream_s2mPipe_ready) begin
        pixelsStream_rValid <= 1'b0;
      end
      if(pixelsStream_s2mPipe_ready) begin
        pixelsStream_s2mPipe_rValid <= pixelsStream_s2mPipe_valid;
      end
      if(when_SuperResolutionPart2_l761) begin
        if(when_SuperResolutionPart2_l763) begin
          outReachRowEnd <= 1'b1;
        end
        if(when_SuperResolutionPart2_l764) begin
          outReachFinalRow <= 1'b1;
        end
        if(when_SuperResolutionPart2_l766) begin
          if(outReachFinalRow) begin
            startRead <= 1'b0;
            readDone <= 1'b1;
            outReachRowEnd <= 1'b0;
            outReachFinalRow <= 1'b0;
          end else begin
            outReachRowEnd <= 1'b0;
          end
        end
        if(controlStream_fire_7) begin
          if(outReachRowEnd) begin
            outReachRowEnd <= 1'b0;
            if(when_SuperResolutionPart2_l783) begin
              oneInFourOutRow <= 1'b1;
            end else begin
              oneInFourOutRow <= 1'b0;
            end
            if(when_SuperResolutionPart2_l785) begin
              twoInFourOutRow <= 1'b1;
            end else begin
              twoInFourOutRow <= 1'b0;
            end
            if(when_SuperResolutionPart2_l787) begin
              threeInFourOutRow <= 1'b1;
            end else begin
              threeInFourOutRow <= 1'b0;
            end
            if(when_SuperResolutionPart2_l789) begin
              zeroInFourOutRow <= 1'b1;
            end else begin
              zeroInFourOutRow <= 1'b0;
            end
          end
          if(when_SuperResolutionPart2_l793) begin
            oneInFourOutPixelAddr <= 1'b1;
          end
          if(oneInFourOutPixelAddr) begin
            oneInFourOutPixelAddr <= 1'b0;
          end
          if(when_SuperResolutionPart2_l796) begin
            twoInFourOutPixelAddr <= 1'b1;
          end
          if(twoInFourOutPixelAddr) begin
            twoInFourOutPixelAddr <= 1'b0;
          end
          if(when_SuperResolutionPart2_l799) begin
            threeInFourOutPixelAddr <= 1'b1;
          end
          if(threeInFourOutPixelAddr) begin
            threeInFourOutPixelAddr <= 1'b0;
          end
          if(when_SuperResolutionPart2_l802) begin
            zeroInFourOutPixelAddr <= 1'b1;
          end
          if(zeroInFourOutPixelAddr) begin
            zeroInFourOutPixelAddr <= 1'b0;
          end
        end
      end
      controlStateMachine_stateReg <= controlStateMachine_stateNext;
      case(controlStateMachine_stateReg)
        controlStateMachine_enumDef_1_HOLD : begin
          if(zeroInFourOutRow) begin
            if(passPixels_fire_13) begin
              if(!threeInFourOutPixelAddr) begin
                holdWillPassToHoldCaseTwo <= 1'b1;
              end
            end
          end else begin
            if(!twoInFourOutRow) begin
              if(threeInFourOutRow) begin
                if(passPixels_fire_15) begin
                  if(threeInFourOutPixelAddr) begin
                    if(willHoldToTwice) begin
                      willHoldToTwice <= 1'b0;
                    end
                  end
                end
              end
            end
          end
          if(passPixels_fire_16) begin
            if(when_SuperResolutionPart2_l560) begin
              willHoldToTwice <= 1'b1;
            end else begin
              willHoldToTwice <= 1'b0;
            end
          end
        end
        controlStateMachine_enumDef_1_PASS : begin
          if(controlStream_fire_8) begin
            if(!oneInFourOutPixelAddr) begin
              if(twoInFourOutPixelAddr) begin
                if(oneInFourOutRow) begin
                  if(when_SuperResolutionPart2_l585) begin
                    willOnceToHoldCaseOne <= 1'b1;
                  end
                end else begin
                  if(twoInFourOutRow) begin
                    if(when_SuperResolutionPart2_l588) begin
                      willOnceToHoldCaseTwo <= 1'b1;
                    end
                  end else begin
                    if(when_SuperResolutionPart2_l590) begin
                      holdWillPassToHoldCaseTwo <= 1'b0;
                    end
                  end
                end
              end
            end
            willPassToHoldCaseOne <= 1'b0;
            willPassToHoldCaseTwo <= 1'b0;
          end
          if(when_SuperResolutionPart2_l602) begin
            willPassToHoldCaseOne <= 1'b1;
          end
          if(when_SuperResolutionPart2_l603) begin
            willPassToHoldCaseOne <= 1'b1;
          end
          if(when_SuperResolutionPart2_l605) begin
            willPassToHoldCaseTwo <= 1'b1;
          end
          if(when_SuperResolutionPart2_l606) begin
            willPassToHoldCaseTwo <= 1'b1;
          end
          if(when_SuperResolutionPart2_l630) begin
            frameStart <= 1'b0;
          end
        end
        controlStateMachine_enumDef_1_ONCE : begin
          if(controlStream_fire_10) begin
            willOnceToHoldCaseOne <= 1'b0;
            willOnceToHoldCaseTwo <= 1'b0;
            willOnceToHoldCaseThree <= 1'b0;
          end
          if(when_SuperResolutionPart2_l662) begin
            willOnceToHoldCaseOne <= 1'b0;
            willOnceToHoldCaseTwo <= 1'b0;
          end
          if(when_SuperResolutionPart2_l667) begin
            willOnceToHoldCaseThree <= 1'b1;
          end
          if(when_SuperResolutionPart2_l668) begin
            willOnceToHoldCaseThree <= 1'b1;
          end
        end
        controlStateMachine_enumDef_1_TWICE : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(posedge clk) begin
    startIn_regNext <= startIn;
    startIn_regNext_1 <= startIn;
    startIn_regNext_2 <= startIn;
    startIn_regNext_3 <= startIn;
    startIn_regNext_4 <= startIn;
    startIn_regNext_5 <= startIn;
    startIn_regNext_6 <= startIn;
    startIn_regNext_7 <= startIn;
    startIn_regNext_8 <= startIn;
    startIn_regNext_9 <= startIn;
    startIn_regNext_10 <= startIn;
    startIn_regNext_11 <= startIn;
    startIn_regNext_12 <= startIn;
    startIn_regNext_13 <= startIn;
    startIn_regNext_14 <= startIn;
    startIn_regNext_15 <= startIn;
    startIn_regNext_16 <= startIn;
    if(pixelsIn_ready) begin
      pixelsIn_rData_pixel <= pixelsIn_payload_pixel;
      pixelsIn_rData_frameStart <= pixelsIn_payload_frameStart;
      pixelsIn_rData_rowEnd <= pixelsIn_payload_rowEnd;
    end
    if(pixelsIn_s2mPipe_ready) begin
      pixelsIn_s2mPipe_rData_pixel <= pixelsIn_s2mPipe_payload_pixel;
      pixelsIn_s2mPipe_rData_frameStart <= pixelsIn_s2mPipe_payload_frameStart;
      pixelsIn_s2mPipe_rData_rowEnd <= pixelsIn_s2mPipe_payload_rowEnd;
    end
    if(mainAddrOneStream_ready) begin
      mainAddrOneStream_rData <= mainAddrOneStream_payload;
    end
    if(mainAddrOneStream_s2mPipe_ready) begin
      mainAddrOneStream_s2mPipe_rData <= mainAddrOneStream_s2mPipe_payload;
    end
    if(CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_mainOnePixelStream_payload_1 <= CICC1851_readStage_mainOnePixelStream_payload;
    end
    if(CICC1851_1) begin
      CICC1851_readStage_mainOnePixelStream_payload_2 <= (CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_mainOnePixelStream_payload_1 : CICC1851_readStage_mainOnePixelStream_payload);
    end
    if(counterAddrOneStream_ready) begin
      counterAddrOneStream_rData <= counterAddrOneStream_payload;
    end
    if(counterAddrOneStream_s2mPipe_ready) begin
      counterAddrOneStream_s2mPipe_rData <= counterAddrOneStream_s2mPipe_payload;
    end
    if(CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_counterOnePixelStream_payload_1 <= CICC1851_readStage_counterOnePixelStream_payload;
    end
    if(CICC1851_2) begin
      CICC1851_readStage_counterOnePixelStream_payload_2 <= (CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_counterOnePixelStream_payload_1 : CICC1851_readStage_counterOnePixelStream_payload);
    end
    if(mainAddrTwoStream_ready) begin
      mainAddrTwoStream_rData <= mainAddrTwoStream_payload;
    end
    if(mainAddrTwoStream_s2mPipe_ready) begin
      mainAddrTwoStream_s2mPipe_rData <= mainAddrTwoStream_s2mPipe_payload;
    end
    if(CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_mainTwoPixelStream_payload_1 <= CICC1851_readStage_mainTwoPixelStream_payload;
    end
    if(CICC1851_3) begin
      CICC1851_readStage_mainTwoPixelStream_payload_2 <= (CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_mainTwoPixelStream_payload_1 : CICC1851_readStage_mainTwoPixelStream_payload);
    end
    if(counterAddrTwoStream_ready) begin
      counterAddrTwoStream_rData <= counterAddrTwoStream_payload;
    end
    if(counterAddrTwoStream_s2mPipe_ready) begin
      counterAddrTwoStream_s2mPipe_rData <= counterAddrTwoStream_s2mPipe_payload;
    end
    if(CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_counterTwoPixelStream_payload_1 <= CICC1851_readStage_counterTwoPixelStream_payload;
    end
    if(CICC1851_4) begin
      CICC1851_readStage_counterTwoPixelStream_payload_2 <= (CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_counterTwoPixelStream_payload_1 : CICC1851_readStage_counterTwoPixelStream_payload);
    end
    if(oddAddrStream_ready) begin
      oddAddrStream_rData <= oddAddrStream_payload;
    end
    if(oddAddrStream_s2mPipe_ready) begin
      oddAddrStream_s2mPipe_rData <= oddAddrStream_s2mPipe_payload;
    end
    if(CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_oddRowPixelStream_payload_1 <= CICC1851_readStage_oddRowPixelStream_payload;
    end
    if(CICC1851_5) begin
      CICC1851_readStage_oddRowPixelStream_payload_2 <= (CICC1851_oddAddrStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_oddRowPixelStream_payload_1 : CICC1851_readStage_oddRowPixelStream_payload);
    end
    if(controlStream_ready) begin
      controlStream_rData_frameStart <= controlStream_payload_frameStart;
      controlStream_rData_rowEnd <= controlStream_payload_rowEnd;
      controlStream_rData_passMode <= controlStream_payload_passMode;
      controlStream_rData_passValid <= controlStream_payload_passValid;
      controlStream_rData_onceMode <= controlStream_payload_onceMode;
      controlStream_rData_onceValid <= controlStream_payload_onceValid;
      controlStream_rData_mainCompare <= controlStream_payload_mainCompare;
      controlStream_rData_counterCompare <= controlStream_payload_counterCompare;
      controlStream_rData_mainDiff <= controlStream_payload_mainDiff;
      controlStream_rData_counterDiff <= controlStream_payload_counterDiff;
      controlStream_rData_twiceCompValid <= controlStream_payload_twiceCompValid;
      controlStream_rData_twiceMode <= controlStream_payload_twiceMode;
      controlStream_rData_inpValidFlag <= controlStream_payload_inpValidFlag;
      controlStream_rData_oddValid <= controlStream_payload_oddValid;
    end
    if(controlStream_s2mPipe_ready) begin
      controlStream_s2mPipe_rData_frameStart <= controlStream_s2mPipe_payload_frameStart;
      controlStream_s2mPipe_rData_rowEnd <= controlStream_s2mPipe_payload_rowEnd;
      controlStream_s2mPipe_rData_passMode <= controlStream_s2mPipe_payload_passMode;
      controlStream_s2mPipe_rData_passValid <= controlStream_s2mPipe_payload_passValid;
      controlStream_s2mPipe_rData_onceMode <= controlStream_s2mPipe_payload_onceMode;
      controlStream_s2mPipe_rData_onceValid <= controlStream_s2mPipe_payload_onceValid;
      controlStream_s2mPipe_rData_mainCompare <= controlStream_s2mPipe_payload_mainCompare;
      controlStream_s2mPipe_rData_counterCompare <= controlStream_s2mPipe_payload_counterCompare;
      controlStream_s2mPipe_rData_mainDiff <= controlStream_s2mPipe_payload_mainDiff;
      controlStream_s2mPipe_rData_counterDiff <= controlStream_s2mPipe_payload_counterDiff;
      controlStream_s2mPipe_rData_twiceCompValid <= controlStream_s2mPipe_payload_twiceCompValid;
      controlStream_s2mPipe_rData_twiceMode <= controlStream_s2mPipe_payload_twiceMode;
      controlStream_s2mPipe_rData_inpValidFlag <= controlStream_s2mPipe_payload_inpValidFlag;
      controlStream_s2mPipe_rData_oddValid <= controlStream_s2mPipe_payload_oddValid;
    end
    if(controlStream_s2mPipe_m2sPipe_ready) begin
      controlStream_s2mPipe_m2sPipe_rData_frameStart <= controlStream_s2mPipe_m2sPipe_payload_frameStart;
      controlStream_s2mPipe_m2sPipe_rData_rowEnd <= controlStream_s2mPipe_m2sPipe_payload_rowEnd;
      controlStream_s2mPipe_m2sPipe_rData_passMode <= controlStream_s2mPipe_m2sPipe_payload_passMode;
      controlStream_s2mPipe_m2sPipe_rData_passValid <= controlStream_s2mPipe_m2sPipe_payload_passValid;
      controlStream_s2mPipe_m2sPipe_rData_onceMode <= controlStream_s2mPipe_m2sPipe_payload_onceMode;
      controlStream_s2mPipe_m2sPipe_rData_onceValid <= controlStream_s2mPipe_m2sPipe_payload_onceValid;
      controlStream_s2mPipe_m2sPipe_rData_mainCompare <= controlStream_s2mPipe_m2sPipe_payload_mainCompare;
      controlStream_s2mPipe_m2sPipe_rData_counterCompare <= controlStream_s2mPipe_m2sPipe_payload_counterCompare;
      controlStream_s2mPipe_m2sPipe_rData_mainDiff <= controlStream_s2mPipe_m2sPipe_payload_mainDiff;
      controlStream_s2mPipe_m2sPipe_rData_counterDiff <= controlStream_s2mPipe_m2sPipe_payload_counterDiff;
      controlStream_s2mPipe_m2sPipe_rData_twiceCompValid <= controlStream_s2mPipe_m2sPipe_payload_twiceCompValid;
      controlStream_s2mPipe_m2sPipe_rData_twiceMode <= controlStream_s2mPipe_m2sPipe_payload_twiceMode;
      controlStream_s2mPipe_m2sPipe_rData_inpValidFlag <= controlStream_s2mPipe_m2sPipe_payload_inpValidFlag;
      controlStream_s2mPipe_m2sPipe_rData_oddValid <= controlStream_s2mPipe_m2sPipe_payload_oddValid;
    end
    if(controlStream_s2mPipe_m2sPipe_m2sPipe_ready) begin
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_frameStart <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_frameStart;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_rowEnd <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_rowEnd;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_passMode <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passMode;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_passValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_onceMode <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceMode;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_onceValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_twiceCompValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceCompValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_twiceMode <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceMode;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_inpValidFlag <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_inpValidFlag;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_oddValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_oddValid;
    end
    if(controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready) begin
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_frameStart <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_frameStart;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_rowEnd <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_rowEnd;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_passMode <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_passMode;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_passValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_passValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_onceMode <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_onceMode;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_onceValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_onceValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_twiceCompValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_twiceCompValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_twiceMode <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_twiceMode;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_inpValidFlag <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_inpValidFlag;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_oddValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_oddValid;
    end
    if(readStage_mainOnePixelStream_ready) begin
      readStage_mainOnePixelStream_rData <= readStage_mainOnePixelStream_payload;
    end
    if(readStage_mainOnePixelStream_s2mPipe_ready) begin
      readStage_mainOnePixelStream_s2mPipe_rData <= readStage_mainOnePixelStream_s2mPipe_payload;
    end
    if(readStage_counterOnePixelStream_ready) begin
      readStage_counterOnePixelStream_rData <= readStage_counterOnePixelStream_payload;
    end
    if(readStage_counterOnePixelStream_s2mPipe_ready) begin
      readStage_counterOnePixelStream_s2mPipe_rData <= readStage_counterOnePixelStream_s2mPipe_payload;
    end
    if(readStage_mainTwoPixelStream_ready) begin
      readStage_mainTwoPixelStream_rData <= readStage_mainTwoPixelStream_payload;
    end
    if(readStage_mainTwoPixelStream_s2mPipe_ready) begin
      readStage_mainTwoPixelStream_s2mPipe_rData <= readStage_mainTwoPixelStream_s2mPipe_payload;
    end
    if(readStage_counterTwoPixelStream_ready) begin
      readStage_counterTwoPixelStream_rData <= readStage_counterTwoPixelStream_payload;
    end
    if(readStage_counterTwoPixelStream_s2mPipe_ready) begin
      readStage_counterTwoPixelStream_s2mPipe_rData <= readStage_counterTwoPixelStream_s2mPipe_payload;
    end
    if(readStage_oddRowPixelStream_ready) begin
      readStage_oddRowPixelStream_rData <= readStage_oddRowPixelStream_payload;
    end
    if(readStage_oddRowPixelStream_s2mPipe_ready) begin
      readStage_oddRowPixelStream_s2mPipe_rData <= readStage_oddRowPixelStream_s2mPipe_payload;
    end
    if(readStage_controlPipe_translated_ready) begin
      readStage_controlPipe_translated_rData_frameStart <= readStage_controlPipe_translated_payload_frameStart;
      readStage_controlPipe_translated_rData_rowEnd <= readStage_controlPipe_translated_payload_rowEnd;
      readStage_controlPipe_translated_rData_passMode <= readStage_controlPipe_translated_payload_passMode;
      readStage_controlPipe_translated_rData_passValid <= readStage_controlPipe_translated_payload_passValid;
      readStage_controlPipe_translated_rData_onceMode <= readStage_controlPipe_translated_payload_onceMode;
      readStage_controlPipe_translated_rData_onceValid <= readStage_controlPipe_translated_payload_onceValid;
      readStage_controlPipe_translated_rData_mainCompare <= readStage_controlPipe_translated_payload_mainCompare;
      readStage_controlPipe_translated_rData_counterCompare <= readStage_controlPipe_translated_payload_counterCompare;
      readStage_controlPipe_translated_rData_mainDiff <= readStage_controlPipe_translated_payload_mainDiff;
      readStage_controlPipe_translated_rData_counterDiff <= readStage_controlPipe_translated_payload_counterDiff;
      readStage_controlPipe_translated_rData_twiceCompValid <= readStage_controlPipe_translated_payload_twiceCompValid;
      readStage_controlPipe_translated_rData_twiceMode <= readStage_controlPipe_translated_payload_twiceMode;
      readStage_controlPipe_translated_rData_inpValidFlag <= readStage_controlPipe_translated_payload_inpValidFlag;
      readStage_controlPipe_translated_rData_oddValid <= readStage_controlPipe_translated_payload_oddValid;
    end
    if(readStage_controlPipe_translated_s2mPipe_ready) begin
      readStage_controlPipe_translated_s2mPipe_rData_frameStart <= readStage_controlPipe_translated_s2mPipe_payload_frameStart;
      readStage_controlPipe_translated_s2mPipe_rData_rowEnd <= readStage_controlPipe_translated_s2mPipe_payload_rowEnd;
      readStage_controlPipe_translated_s2mPipe_rData_passMode <= readStage_controlPipe_translated_s2mPipe_payload_passMode;
      readStage_controlPipe_translated_s2mPipe_rData_passValid <= readStage_controlPipe_translated_s2mPipe_payload_passValid;
      readStage_controlPipe_translated_s2mPipe_rData_onceMode <= readStage_controlPipe_translated_s2mPipe_payload_onceMode;
      readStage_controlPipe_translated_s2mPipe_rData_onceValid <= readStage_controlPipe_translated_s2mPipe_payload_onceValid;
      readStage_controlPipe_translated_s2mPipe_rData_mainCompare <= readStage_controlPipe_translated_s2mPipe_payload_mainCompare;
      readStage_controlPipe_translated_s2mPipe_rData_counterCompare <= readStage_controlPipe_translated_s2mPipe_payload_counterCompare;
      readStage_controlPipe_translated_s2mPipe_rData_mainDiff <= readStage_controlPipe_translated_s2mPipe_payload_mainDiff;
      readStage_controlPipe_translated_s2mPipe_rData_counterDiff <= readStage_controlPipe_translated_s2mPipe_payload_counterDiff;
      readStage_controlPipe_translated_s2mPipe_rData_twiceCompValid <= readStage_controlPipe_translated_s2mPipe_payload_twiceCompValid;
      readStage_controlPipe_translated_s2mPipe_rData_twiceMode <= readStage_controlPipe_translated_s2mPipe_payload_twiceMode;
      readStage_controlPipe_translated_s2mPipe_rData_inpValidFlag <= readStage_controlPipe_translated_s2mPipe_payload_inpValidFlag;
      readStage_controlPipe_translated_s2mPipe_rData_oddValid <= readStage_controlPipe_translated_s2mPipe_payload_oddValid;
    end
    if(compareStage_mainOnePixelStream_ready) begin
      compareStage_mainOnePixelStream_rData <= compareStage_mainOnePixelStream_payload;
    end
    if(compareStage_mainOnePixelStream_s2mPipe_ready) begin
      compareStage_mainOnePixelStream_s2mPipe_rData <= compareStage_mainOnePixelStream_s2mPipe_payload;
    end
    if(compareStage_counterOnePixelStream_ready) begin
      compareStage_counterOnePixelStream_rData <= compareStage_counterOnePixelStream_payload;
    end
    if(compareStage_counterOnePixelStream_s2mPipe_ready) begin
      compareStage_counterOnePixelStream_s2mPipe_rData <= compareStage_counterOnePixelStream_s2mPipe_payload;
    end
    if(compareStage_mainTwoPixelStream_ready) begin
      compareStage_mainTwoPixelStream_rData <= compareStage_mainTwoPixelStream_payload;
    end
    if(compareStage_mainTwoPixelStream_s2mPipe_ready) begin
      compareStage_mainTwoPixelStream_s2mPipe_rData <= compareStage_mainTwoPixelStream_s2mPipe_payload;
    end
    if(compareStage_counterTwoPixelStream_ready) begin
      compareStage_counterTwoPixelStream_rData <= compareStage_counterTwoPixelStream_payload;
    end
    if(compareStage_counterTwoPixelStream_s2mPipe_ready) begin
      compareStage_counterTwoPixelStream_s2mPipe_rData <= compareStage_counterTwoPixelStream_s2mPipe_payload;
    end
    if(compareStage_oddRowPixelStream_ready) begin
      compareStage_oddRowPixelStream_rData <= compareStage_oddRowPixelStream_payload;
    end
    if(compareStage_oddRowPixelStream_s2mPipe_ready) begin
      compareStage_oddRowPixelStream_s2mPipe_rData <= compareStage_oddRowPixelStream_s2mPipe_payload;
    end
    if(compareStage_controlPipe_translated_ready) begin
      compareStage_controlPipe_translated_rData_frameStart <= compareStage_controlPipe_translated_payload_frameStart;
      compareStage_controlPipe_translated_rData_rowEnd <= compareStage_controlPipe_translated_payload_rowEnd;
      compareStage_controlPipe_translated_rData_passMode <= compareStage_controlPipe_translated_payload_passMode;
      compareStage_controlPipe_translated_rData_passValid <= compareStage_controlPipe_translated_payload_passValid;
      compareStage_controlPipe_translated_rData_onceMode <= compareStage_controlPipe_translated_payload_onceMode;
      compareStage_controlPipe_translated_rData_onceValid <= compareStage_controlPipe_translated_payload_onceValid;
      compareStage_controlPipe_translated_rData_mainCompare <= compareStage_controlPipe_translated_payload_mainCompare;
      compareStage_controlPipe_translated_rData_counterCompare <= compareStage_controlPipe_translated_payload_counterCompare;
      compareStage_controlPipe_translated_rData_mainDiff <= compareStage_controlPipe_translated_payload_mainDiff;
      compareStage_controlPipe_translated_rData_counterDiff <= compareStage_controlPipe_translated_payload_counterDiff;
      compareStage_controlPipe_translated_rData_twiceCompValid <= compareStage_controlPipe_translated_payload_twiceCompValid;
      compareStage_controlPipe_translated_rData_twiceMode <= compareStage_controlPipe_translated_payload_twiceMode;
      compareStage_controlPipe_translated_rData_inpValidFlag <= compareStage_controlPipe_translated_payload_inpValidFlag;
      compareStage_controlPipe_translated_rData_oddValid <= compareStage_controlPipe_translated_payload_oddValid;
    end
    if(compareStage_controlPipe_translated_s2mPipe_ready) begin
      compareStage_controlPipe_translated_s2mPipe_rData_frameStart <= compareStage_controlPipe_translated_s2mPipe_payload_frameStart;
      compareStage_controlPipe_translated_s2mPipe_rData_rowEnd <= compareStage_controlPipe_translated_s2mPipe_payload_rowEnd;
      compareStage_controlPipe_translated_s2mPipe_rData_passMode <= compareStage_controlPipe_translated_s2mPipe_payload_passMode;
      compareStage_controlPipe_translated_s2mPipe_rData_passValid <= compareStage_controlPipe_translated_s2mPipe_payload_passValid;
      compareStage_controlPipe_translated_s2mPipe_rData_onceMode <= compareStage_controlPipe_translated_s2mPipe_payload_onceMode;
      compareStage_controlPipe_translated_s2mPipe_rData_onceValid <= compareStage_controlPipe_translated_s2mPipe_payload_onceValid;
      compareStage_controlPipe_translated_s2mPipe_rData_mainCompare <= compareStage_controlPipe_translated_s2mPipe_payload_mainCompare;
      compareStage_controlPipe_translated_s2mPipe_rData_counterCompare <= compareStage_controlPipe_translated_s2mPipe_payload_counterCompare;
      compareStage_controlPipe_translated_s2mPipe_rData_mainDiff <= compareStage_controlPipe_translated_s2mPipe_payload_mainDiff;
      compareStage_controlPipe_translated_s2mPipe_rData_counterDiff <= compareStage_controlPipe_translated_s2mPipe_payload_counterDiff;
      compareStage_controlPipe_translated_s2mPipe_rData_twiceCompValid <= compareStage_controlPipe_translated_s2mPipe_payload_twiceCompValid;
      compareStage_controlPipe_translated_s2mPipe_rData_twiceMode <= compareStage_controlPipe_translated_s2mPipe_payload_twiceMode;
      compareStage_controlPipe_translated_s2mPipe_rData_inpValidFlag <= compareStage_controlPipe_translated_s2mPipe_payload_inpValidFlag;
      compareStage_controlPipe_translated_s2mPipe_rData_oddValid <= compareStage_controlPipe_translated_s2mPipe_payload_oddValid;
    end
    if(diffStage_mainOnePixelStream_ready) begin
      diffStage_mainOnePixelStream_rData <= diffStage_mainOnePixelStream_payload;
    end
    if(diffStage_mainOnePixelStream_s2mPipe_ready) begin
      diffStage_mainOnePixelStream_s2mPipe_rData <= diffStage_mainOnePixelStream_s2mPipe_payload;
    end
    if(diffStage_counterOnePixelStream_ready) begin
      diffStage_counterOnePixelStream_rData <= diffStage_counterOnePixelStream_payload;
    end
    if(diffStage_counterOnePixelStream_s2mPipe_ready) begin
      diffStage_counterOnePixelStream_s2mPipe_rData <= diffStage_counterOnePixelStream_s2mPipe_payload;
    end
    if(diffStage_mainTwoPixelStream_ready) begin
      diffStage_mainTwoPixelStream_rData <= diffStage_mainTwoPixelStream_payload;
    end
    if(diffStage_mainTwoPixelStream_s2mPipe_ready) begin
      diffStage_mainTwoPixelStream_s2mPipe_rData <= diffStage_mainTwoPixelStream_s2mPipe_payload;
    end
    if(diffStage_counterTwoPixelStream_ready) begin
      diffStage_counterTwoPixelStream_rData <= diffStage_counterTwoPixelStream_payload;
    end
    if(diffStage_counterTwoPixelStream_s2mPipe_ready) begin
      diffStage_counterTwoPixelStream_s2mPipe_rData <= diffStage_counterTwoPixelStream_s2mPipe_payload;
    end
    if(diffStage_oddRowPixelStream_ready) begin
      diffStage_oddRowPixelStream_rData <= diffStage_oddRowPixelStream_payload;
    end
    if(diffStage_oddRowPixelStream_s2mPipe_ready) begin
      diffStage_oddRowPixelStream_s2mPipe_rData <= diffStage_oddRowPixelStream_s2mPipe_payload;
    end
    if(diffStage_controlPipe_fork_io_outputs_0_translated_ready) begin
      diffStage_controlPipe_fork_io_outputs_0_translated_rData_frameStart <= diffStage_controlPipe_fork_io_outputs_0_translated_payload_frameStart;
      diffStage_controlPipe_fork_io_outputs_0_translated_rData_rowEnd <= diffStage_controlPipe_fork_io_outputs_0_translated_payload_rowEnd;
      diffStage_controlPipe_fork_io_outputs_0_translated_rData_passMode <= diffStage_controlPipe_fork_io_outputs_0_translated_payload_passMode;
      diffStage_controlPipe_fork_io_outputs_0_translated_rData_passValid <= diffStage_controlPipe_fork_io_outputs_0_translated_payload_passValid;
      diffStage_controlPipe_fork_io_outputs_0_translated_rData_onceMode <= diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceMode;
      diffStage_controlPipe_fork_io_outputs_0_translated_rData_onceValid <= diffStage_controlPipe_fork_io_outputs_0_translated_payload_onceValid;
      diffStage_controlPipe_fork_io_outputs_0_translated_rData_mainCompare <= diffStage_controlPipe_fork_io_outputs_0_translated_payload_mainCompare;
      diffStage_controlPipe_fork_io_outputs_0_translated_rData_counterCompare <= diffStage_controlPipe_fork_io_outputs_0_translated_payload_counterCompare;
      diffStage_controlPipe_fork_io_outputs_0_translated_rData_mainDiff <= diffStage_controlPipe_fork_io_outputs_0_translated_payload_mainDiff;
      diffStage_controlPipe_fork_io_outputs_0_translated_rData_counterDiff <= diffStage_controlPipe_fork_io_outputs_0_translated_payload_counterDiff;
      diffStage_controlPipe_fork_io_outputs_0_translated_rData_twiceCompValid <= diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceCompValid;
      diffStage_controlPipe_fork_io_outputs_0_translated_rData_twiceMode <= diffStage_controlPipe_fork_io_outputs_0_translated_payload_twiceMode;
      diffStage_controlPipe_fork_io_outputs_0_translated_rData_inpValidFlag <= diffStage_controlPipe_fork_io_outputs_0_translated_payload_inpValidFlag;
      diffStage_controlPipe_fork_io_outputs_0_translated_rData_oddValid <= diffStage_controlPipe_fork_io_outputs_0_translated_payload_oddValid;
    end
    if(diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_ready) begin
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_frameStart <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_frameStart;
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_rowEnd <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_rowEnd;
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_passMode <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_passMode;
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_passValid <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_passValid;
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_onceMode <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_onceMode;
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_onceValid <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_onceValid;
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_mainCompare <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_mainCompare;
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_counterCompare <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_counterCompare;
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_mainDiff <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_mainDiff;
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_counterDiff <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_counterDiff;
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_twiceCompValid <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_twiceCompValid;
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_twiceMode <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_twiceMode;
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_inpValidFlag <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_inpValidFlag;
      diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_rData_oddValid <= diffStage_controlPipe_fork_io_outputs_0_translated_s2mPipe_payload_oddValid;
    end
    if(resultStage_pixelStream_ready) begin
      resultStage_pixelStream_rData <= resultStage_pixelStream_payload;
    end
    if(resultStage_pixelStream_s2mPipe_ready) begin
      resultStage_pixelStream_s2mPipe_rData <= resultStage_pixelStream_s2mPipe_payload;
    end
    if(pixelsStream_ready) begin
      pixelsStream_rData_pixel <= pixelsStream_payload_pixel;
      pixelsStream_rData_frameStart <= pixelsStream_payload_frameStart;
      pixelsStream_rData_rowEnd <= pixelsStream_payload_rowEnd;
      pixelsStream_rData_inpValid <= pixelsStream_payload_inpValid;
    end
    if(pixelsStream_s2mPipe_ready) begin
      pixelsStream_s2mPipe_rData_pixel <= pixelsStream_s2mPipe_payload_pixel;
      pixelsStream_s2mPipe_rData_frameStart <= pixelsStream_s2mPipe_payload_frameStart;
      pixelsStream_s2mPipe_rData_rowEnd <= pixelsStream_s2mPipe_payload_rowEnd;
      pixelsStream_s2mPipe_rData_inpValid <= pixelsStream_s2mPipe_payload_inpValid;
    end
  end


endmodule

module SuperResolutionPart1 (
  input               pixelsIn_valid,
  output reg          pixelsIn_ready,
  input      [7:0]    pixelsIn_payload_pixel,
  input               pixelsIn_payload_frameStart,
  input               pixelsIn_payload_rowEnd,
  input               startIn,
  input               inpTwoDoneIn,
  input               inpThreeDoneIn,
  output reg          pixelsOut_valid,
  input               pixelsOut_ready,
  output reg [7:0]    pixelsOut_payload_pixel,
  output reg          pixelsOut_payload_frameStart,
  output reg          pixelsOut_payload_rowEnd,
  output reg          startOut,
  output reg          inpDoneOut,
  input      [7:0]    thresholdIn,
  input      [9:0]    widthIn,
  input      [9:0]    heightIn,
  input               clk,
  input               resetn
);
  localparam controlStateMachine_enumDef_BOOT = 3'd0;
  localparam controlStateMachine_enumDef_HOLD = 3'd1;
  localparam controlStateMachine_enumDef_PASS = 3'd2;
  localparam controlStateMachine_enumDef_ONCE = 3'd3;
  localparam controlStateMachine_enumDef_TWICE = 3'd4;

  wire                diffStage_controlPipe_fork_io_outputs_0_ready;
  reg        [7:0]    CICC1851_lineBufferOne_port0;
  reg        [7:0]    CICC1851_lineBufferOne_port1;
  reg        [7:0]    CICC1851_lineBufferTwo_port0;
  reg        [7:0]    CICC1851_lineBufferTwo_port1;
  wire                diffStage_controlPipe_fork_io_input_ready;
  wire                diffStage_controlPipe_fork_io_outputs_0_valid;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_frameStart;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_rowEnd;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_passMode;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_passValid;
  wire       [2:0]    diffStage_controlPipe_fork_io_outputs_0_payload_onceMode;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_onceValid;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_mainCompare;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_counterCompare;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_payload_mainDiff;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_payload_counterDiff;
  wire                diffStage_controlPipe_fork_io_outputs_0_payload_twiceCompValid;
  wire       [2:0]    diffStage_controlPipe_fork_io_outputs_0_payload_twiceMode;
  wire                diffStage_controlPipe_fork_io_outputs_1_valid;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_frameStart;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_rowEnd;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_passMode;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_passValid;
  wire       [2:0]    diffStage_controlPipe_fork_io_outputs_1_payload_onceMode;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_onceValid;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_mainCompare;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_counterCompare;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff;
  wire                diffStage_controlPipe_fork_io_outputs_1_payload_twiceCompValid;
  wire       [2:0]    diffStage_controlPipe_fork_io_outputs_1_payload_twiceMode;
  wire       [9:0]    CICC1851_bufferRowCount_valueNext;
  wire       [0:0]    CICC1851_bufferRowCount_valueNext_1;
  wire       [9:0]    CICC1851_bufferWAddr_valueNext;
  wire       [0:0]    CICC1851_bufferWAddr_valueNext_1;
  wire       [10:0]   CICC1851_outPixelAddr_valueNext;
  wire       [0:0]    CICC1851_outPixelAddr_valueNext_1;
  wire       [10:0]   CICC1851_outRowCount_valueNext;
  wire       [0:0]    CICC1851_outRowCount_valueNext_1;
  wire       [10:0]   CICC1851_mainAddrOne;
  wire       [10:0]   CICC1851_counterAddrOne;
  wire       [10:0]   CICC1851_mainAddrTwo;
  wire       [10:0]   CICC1851_counterAddrTwo;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_1;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_2;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_3;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_4;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_5;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_6;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_7;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_8;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_9;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_10;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_11;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_12;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_13;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_14;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_15;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_16;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_17;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_18;
  wire       [8:0]    CICC1851_resultStage_pixelStream_payload_19;
  wire       [9:0]    CICC1851_when_SuperResolutionPart1_l421;
  wire       [9:0]    CICC1851_when_SuperResolutionPart1_l422;
  wire       [10:0]   CICC1851_when_SuperResolutionPart1_l447;
  wire       [7:0]    CICC1851_lineBufferTwo_port;
  wire                CICC1851_lineBufferTwo_port_1;
  wire       [7:0]    CICC1851_lineBufferOne_port;
  wire                CICC1851_lineBufferOne_port_1;
  wire       [10:0]   CICC1851_when_SuperResolutionPart1_l482;
  wire       [10:0]   CICC1851_when_SuperResolutionPart1_l484;
  wire       [10:0]   CICC1851_when_SuperResolutionPart1_l489;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l498;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l498_1;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l500;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l500_1;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l500_2;
  wire       [2:0]    CICC1851_when_SuperResolutionPart1_l500_3;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l510;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l510_1;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l510_2;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l511;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l511_1;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l511_2;
  wire       [10:0]   CICC1851_when_SuperResolutionPart1_l537;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l542;
  wire       [10:0]   CICC1851_when_SuperResolutionPart1_l542_1;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l542_2;
  wire       [10:0]   CICC1851_mainAddrOne_1;
  wire       [10:0]   CICC1851_mainAddrOne_2;
  wire       [10:0]   CICC1851_counterAddrOne_1;
  wire       [10:0]   CICC1851_counterAddrOne_2;
  wire       [11:0]   CICC1851_counterAddrOne_3;
  wire       [11:0]   CICC1851_counterAddrOne_4;
  wire       [11:0]   CICC1851_counterAddrOne_5;
  wire       [1:0]    CICC1851_counterAddrOne_6;
  wire       [0:0]    CICC1851_controls_onceMode;
  wire       [10:0]   CICC1851_mainAddrTwo_1;
  wire       [10:0]   CICC1851_mainAddrTwo_2;
  wire       [10:0]   CICC1851_counterAddrTwo_1;
  wire       [10:0]   CICC1851_counterAddrTwo_2;
  wire       [11:0]   CICC1851_counterAddrTwo_3;
  wire       [11:0]   CICC1851_counterAddrTwo_4;
  wire       [11:0]   CICC1851_counterAddrTwo_5;
  wire       [1:0]    CICC1851_counterAddrTwo_6;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l563;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l563_1;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l563_2;
  wire       [2:0]    CICC1851_when_SuperResolutionPart1_l563_3;
  wire       [1:0]    CICC1851_controls_onceMode_1;
  wire       [1:0]    CICC1851_controls_onceMode_2;
  wire       [10:0]   CICC1851_mainAddrOne_3;
  wire       [10:0]   CICC1851_mainAddrTwo_3;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l578;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l578_1;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l578_2;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l579;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l579_1;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l579_2;
  wire       [10:0]   CICC1851_mainAddrOne_4;
  wire       [10:0]   CICC1851_mainAddrOne_5;
  wire       [10:0]   CICC1851_mainAddrOne_6;
  wire       [10:0]   CICC1851_mainAddrOne_7;
  wire       [11:0]   CICC1851_counterAddrOne_7;
  wire       [11:0]   CICC1851_counterAddrOne_8;
  wire       [11:0]   CICC1851_counterAddrOne_9;
  wire       [1:0]    CICC1851_counterAddrOne_10;
  wire       [10:0]   CICC1851_mainAddrTwo_4;
  wire       [10:0]   CICC1851_mainAddrTwo_5;
  wire       [10:0]   CICC1851_mainAddrTwo_6;
  wire       [10:0]   CICC1851_mainAddrTwo_7;
  wire       [11:0]   CICC1851_counterAddrTwo_7;
  wire       [11:0]   CICC1851_counterAddrTwo_8;
  wire       [11:0]   CICC1851_counterAddrTwo_9;
  wire       [1:0]    CICC1851_counterAddrTwo_10;
  wire       [10:0]   CICC1851_mainAddrOne_8;
  wire       [10:0]   CICC1851_mainAddrOne_9;
  wire       [10:0]   CICC1851_counterAddrTwo_11;
  wire       [10:0]   CICC1851_counterAddrTwo_12;
  wire       [10:0]   CICC1851_mainAddrTwo_8;
  wire       [10:0]   CICC1851_mainAddrTwo_9;
  wire       [10:0]   CICC1851_counterAddrOne_11;
  wire       [10:0]   CICC1851_counterAddrOne_12;
  wire       [11:0]   CICC1851_mainAddrTwo_10;
  wire       [11:0]   CICC1851_mainAddrTwo_11;
  wire       [11:0]   CICC1851_mainAddrTwo_12;
  wire       [1:0]    CICC1851_mainAddrTwo_13;
  wire       [11:0]   CICC1851_counterAddrOne_13;
  wire       [11:0]   CICC1851_counterAddrOne_14;
  wire       [11:0]   CICC1851_counterAddrOne_15;
  wire       [1:0]    CICC1851_counterAddrOne_16;
  wire       [10:0]   CICC1851_mainAddrTwo_14;
  wire       [10:0]   CICC1851_mainAddrTwo_15;
  wire       [10:0]   CICC1851_counterAddrOne_17;
  wire       [10:0]   CICC1851_counterAddrOne_18;
  wire       [10:0]   CICC1851_mainAddrOne_10;
  wire       [10:0]   CICC1851_mainAddrOne_11;
  wire       [10:0]   CICC1851_counterAddrTwo_13;
  wire       [10:0]   CICC1851_counterAddrTwo_14;
  wire       [11:0]   CICC1851_mainAddrOne_12;
  wire       [11:0]   CICC1851_mainAddrOne_13;
  wire       [11:0]   CICC1851_mainAddrOne_14;
  wire       [1:0]    CICC1851_mainAddrOne_15;
  wire       [11:0]   CICC1851_counterAddrTwo_15;
  wire       [11:0]   CICC1851_counterAddrTwo_16;
  wire       [11:0]   CICC1851_counterAddrTwo_17;
  wire       [1:0]    CICC1851_counterAddrTwo_18;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l664;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l664_1;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l664_2;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l665;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l665_1;
  wire       [11:0]   CICC1851_when_SuperResolutionPart1_l665_2;
  reg                 inpDone;
  wire                when_SuperResolutionPart1_l79;
  reg                 startIn_regNext;
  wire                when_SuperResolutionPart1_l79_1;
  reg                 readDone;
  wire                when_SuperResolutionPart1_l82;
  reg                 startRead;
  wire                when_SuperResolutionPart1_l85;
  wire                when_SuperResolutionPart1_l85_1;
  reg                 slaveStart;
  wire                pixelsIn_fire;
  wire                when_SuperResolutionPart1_l88;
  wire                when_SuperResolutionPart1_l88_1;
  reg                 frameStart;
  reg        [7:0]    inpThreshold;
  reg        [9:0]    bmpWidth;
  reg        [9:0]    bmpHeight;
  reg                 holdBuffer;
  wire                when_SuperResolutionPart1_l103;
  reg                 writeDone;
  wire                when_SuperResolutionPart1_l106;
  reg                 bufferRowCount_willIncrement;
  reg                 bufferRowCount_willClear;
  reg        [9:0]    bufferRowCount_valueNext;
  reg        [9:0]    bufferRowCount_value;
  wire                bufferRowCount_willOverflowIfInc;
  wire                bufferRowCount_willOverflow;
  reg                 bufferEnable;
  wire                when_SuperResolutionPart1_l112;
  wire                when_SuperResolutionPart1_l112_1;
  reg                 bufferSwitch;
  wire                when_SuperResolutionPart1_l115;
  reg                 nextRowBuffer;
  wire                when_SuperResolutionPart1_l118;
  reg                 bufferReuse;
  reg                 bufferWAddr_willIncrement;
  reg                 bufferWAddr_willClear;
  reg        [9:0]    bufferWAddr_valueNext;
  reg        [9:0]    bufferWAddr_value;
  wire                bufferWAddr_willOverflowIfInc;
  wire                bufferWAddr_willOverflow;
  reg                 outPixelAddr_willIncrement;
  reg                 outPixelAddr_willClear;
  reg        [10:0]   outPixelAddr_valueNext;
  reg        [10:0]   outPixelAddr_value;
  wire                outPixelAddr_willOverflowIfInc;
  wire                outPixelAddr_willOverflow;
  reg                 outRowCount_willIncrement;
  reg                 outRowCount_willClear;
  reg        [10:0]   outRowCount_valueNext;
  reg        [10:0]   outRowCount_value;
  wire                outRowCount_willOverflowIfInc;
  wire                outRowCount_willOverflow;
  reg                 outReachRowEnd;
  reg                 outReachFinalRow;
  reg                 bufferReachRowEnd;
  reg                 bufferReachFinalRow;
  reg        [9:0]    mainAddrOne;
  reg        [9:0]    counterAddrOne;
  reg        [9:0]    mainAddrTwo;
  reg        [9:0]    counterAddrTwo;
  wire                validStream_valid;
  reg                 validStream_ready;
  wire                controlStream_valid;
  wire                controlStream_ready;
  wire                controlStream_payload_frameStart;
  wire                controlStream_payload_rowEnd;
  wire                controlStream_payload_passMode;
  wire                controlStream_payload_passValid;
  wire       [2:0]    controlStream_payload_onceMode;
  wire                controlStream_payload_onceValid;
  wire                controlStream_payload_mainCompare;
  wire                controlStream_payload_counterCompare;
  wire       [7:0]    controlStream_payload_mainDiff;
  wire       [7:0]    controlStream_payload_counterDiff;
  wire                controlStream_payload_twiceCompValid;
  wire       [2:0]    controlStream_payload_twiceMode;
  reg                 controls_frameStart;
  reg                 controls_rowEnd;
  reg                 controls_passMode;
  reg                 controls_passValid;
  reg        [2:0]    controls_onceMode;
  reg                 controls_onceValid;
  wire                controls_mainCompare;
  wire                controls_counterCompare;
  wire       [7:0]    controls_mainDiff;
  wire       [7:0]    controls_counterDiff;
  reg                 controls_twiceCompValid;
  reg        [2:0]    controls_twiceMode;
  wire       [29:0]   CICC1851_controls_frameStart;
  wire                mainAddrOneStream_valid;
  wire                mainAddrOneStream_ready;
  wire       [9:0]    mainAddrOneStream_payload;
  wire                counterAddrOneStream_valid;
  wire                counterAddrOneStream_ready;
  wire       [9:0]    counterAddrOneStream_payload;
  wire                mainAddrTwoStream_valid;
  wire                mainAddrTwoStream_ready;
  wire       [9:0]    mainAddrTwoStream_payload;
  wire                counterAddrTwoStream_valid;
  wire                counterAddrTwoStream_ready;
  wire       [9:0]    counterAddrTwoStream_payload;
  wire                mainAddrOneStream_s2mPipe_valid;
  reg                 mainAddrOneStream_s2mPipe_ready;
  wire       [9:0]    mainAddrOneStream_s2mPipe_payload;
  reg                 mainAddrOneStream_rValid;
  reg        [9:0]    mainAddrOneStream_rData;
  wire                mainAddrOneStream_s2mPipe_m2sPipe_valid;
  wire                mainAddrOneStream_s2mPipe_m2sPipe_ready;
  wire       [9:0]    mainAddrOneStream_s2mPipe_m2sPipe_payload;
  reg                 mainAddrOneStream_s2mPipe_rValid;
  reg        [9:0]    mainAddrOneStream_s2mPipe_rData;
  wire                when_Stream_l368;
  wire                CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_mainOnePixelStream_payload;
  reg                 CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_1;
  reg                 CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_mainOnePixelStream_payload_1;
  wire                readStage_mainOnePixelStream_valid;
  wire                readStage_mainOnePixelStream_ready;
  wire       [7:0]    readStage_mainOnePixelStream_payload;
  reg                 CICC1851_readStage_mainOnePixelStream_valid;
  reg        [7:0]    CICC1851_readStage_mainOnePixelStream_payload_2;
  wire                when_Stream_l368_1;
  wire                counterAddrOneStream_s2mPipe_valid;
  reg                 counterAddrOneStream_s2mPipe_ready;
  wire       [9:0]    counterAddrOneStream_s2mPipe_payload;
  reg                 counterAddrOneStream_rValid;
  reg        [9:0]    counterAddrOneStream_rData;
  wire                counterAddrOneStream_s2mPipe_m2sPipe_valid;
  wire                counterAddrOneStream_s2mPipe_m2sPipe_ready;
  wire       [9:0]    counterAddrOneStream_s2mPipe_m2sPipe_payload;
  reg                 counterAddrOneStream_s2mPipe_rValid;
  reg        [9:0]    counterAddrOneStream_s2mPipe_rData;
  wire                when_Stream_l368_2;
  wire                CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_counterOnePixelStream_payload;
  reg                 CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_2;
  reg                 CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_counterOnePixelStream_payload_1;
  wire                readStage_counterOnePixelStream_valid;
  wire                readStage_counterOnePixelStream_ready;
  wire       [7:0]    readStage_counterOnePixelStream_payload;
  reg                 CICC1851_readStage_counterOnePixelStream_valid;
  reg        [7:0]    CICC1851_readStage_counterOnePixelStream_payload_2;
  wire                when_Stream_l368_3;
  wire                mainAddrTwoStream_s2mPipe_valid;
  reg                 mainAddrTwoStream_s2mPipe_ready;
  wire       [9:0]    mainAddrTwoStream_s2mPipe_payload;
  reg                 mainAddrTwoStream_rValid;
  reg        [9:0]    mainAddrTwoStream_rData;
  wire                mainAddrTwoStream_s2mPipe_m2sPipe_valid;
  wire                mainAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire       [9:0]    mainAddrTwoStream_s2mPipe_m2sPipe_payload;
  reg                 mainAddrTwoStream_s2mPipe_rValid;
  reg        [9:0]    mainAddrTwoStream_s2mPipe_rData;
  wire                when_Stream_l368_4;
  wire                CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_mainTwoPixelStream_payload;
  reg                 CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_3;
  reg                 CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_mainTwoPixelStream_payload_1;
  wire                readStage_mainTwoPixelStream_valid;
  wire                readStage_mainTwoPixelStream_ready;
  wire       [7:0]    readStage_mainTwoPixelStream_payload;
  reg                 CICC1851_readStage_mainTwoPixelStream_valid;
  reg        [7:0]    CICC1851_readStage_mainTwoPixelStream_payload_2;
  wire                when_Stream_l368_5;
  wire                counterAddrTwoStream_s2mPipe_valid;
  reg                 counterAddrTwoStream_s2mPipe_ready;
  wire       [9:0]    counterAddrTwoStream_s2mPipe_payload;
  reg                 counterAddrTwoStream_rValid;
  reg        [9:0]    counterAddrTwoStream_rData;
  wire                counterAddrTwoStream_s2mPipe_m2sPipe_valid;
  wire                counterAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire       [9:0]    counterAddrTwoStream_s2mPipe_m2sPipe_payload;
  reg                 counterAddrTwoStream_s2mPipe_rValid;
  reg        [9:0]    counterAddrTwoStream_s2mPipe_rData;
  wire                when_Stream_l368_6;
  wire                CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready;
  wire                CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_1;
  wire       [7:0]    CICC1851_readStage_counterTwoPixelStream_payload;
  reg                 CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  reg                 CICC1851_4;
  reg                 CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_3;
  reg        [7:0]    CICC1851_readStage_counterTwoPixelStream_payload_1;
  wire                readStage_counterTwoPixelStream_valid;
  wire                readStage_counterTwoPixelStream_ready;
  wire       [7:0]    readStage_counterTwoPixelStream_payload;
  reg                 CICC1851_readStage_counterTwoPixelStream_valid;
  reg        [7:0]    CICC1851_readStage_counterTwoPixelStream_payload_2;
  wire                when_Stream_l368_7;
  wire                controlStream_s2mPipe_valid;
  reg                 controlStream_s2mPipe_ready;
  wire                controlStream_s2mPipe_payload_frameStart;
  wire                controlStream_s2mPipe_payload_rowEnd;
  wire                controlStream_s2mPipe_payload_passMode;
  wire                controlStream_s2mPipe_payload_passValid;
  wire       [2:0]    controlStream_s2mPipe_payload_onceMode;
  wire                controlStream_s2mPipe_payload_onceValid;
  wire                controlStream_s2mPipe_payload_mainCompare;
  wire                controlStream_s2mPipe_payload_counterCompare;
  wire       [7:0]    controlStream_s2mPipe_payload_mainDiff;
  wire       [7:0]    controlStream_s2mPipe_payload_counterDiff;
  wire                controlStream_s2mPipe_payload_twiceCompValid;
  wire       [2:0]    controlStream_s2mPipe_payload_twiceMode;
  reg                 controlStream_rValid;
  reg                 controlStream_rData_frameStart;
  reg                 controlStream_rData_rowEnd;
  reg                 controlStream_rData_passMode;
  reg                 controlStream_rData_passValid;
  reg        [2:0]    controlStream_rData_onceMode;
  reg                 controlStream_rData_onceValid;
  reg                 controlStream_rData_mainCompare;
  reg                 controlStream_rData_counterCompare;
  reg        [7:0]    controlStream_rData_mainDiff;
  reg        [7:0]    controlStream_rData_counterDiff;
  reg                 controlStream_rData_twiceCompValid;
  reg        [2:0]    controlStream_rData_twiceMode;
  wire                controlStream_s2mPipe_m2sPipe_valid;
  reg                 controlStream_s2mPipe_m2sPipe_ready;
  wire                controlStream_s2mPipe_m2sPipe_payload_frameStart;
  wire                controlStream_s2mPipe_m2sPipe_payload_rowEnd;
  wire                controlStream_s2mPipe_m2sPipe_payload_passMode;
  wire                controlStream_s2mPipe_m2sPipe_payload_passValid;
  wire       [2:0]    controlStream_s2mPipe_m2sPipe_payload_onceMode;
  wire                controlStream_s2mPipe_m2sPipe_payload_onceValid;
  wire                controlStream_s2mPipe_m2sPipe_payload_mainCompare;
  wire                controlStream_s2mPipe_m2sPipe_payload_counterCompare;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_payload_mainDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_payload_counterDiff;
  wire                controlStream_s2mPipe_m2sPipe_payload_twiceCompValid;
  wire       [2:0]    controlStream_s2mPipe_m2sPipe_payload_twiceMode;
  reg                 controlStream_s2mPipe_rValid;
  reg                 controlStream_s2mPipe_rData_frameStart;
  reg                 controlStream_s2mPipe_rData_rowEnd;
  reg                 controlStream_s2mPipe_rData_passMode;
  reg                 controlStream_s2mPipe_rData_passValid;
  reg        [2:0]    controlStream_s2mPipe_rData_onceMode;
  reg                 controlStream_s2mPipe_rData_onceValid;
  reg                 controlStream_s2mPipe_rData_mainCompare;
  reg                 controlStream_s2mPipe_rData_counterCompare;
  reg        [7:0]    controlStream_s2mPipe_rData_mainDiff;
  reg        [7:0]    controlStream_s2mPipe_rData_counterDiff;
  reg                 controlStream_s2mPipe_rData_twiceCompValid;
  reg        [2:0]    controlStream_s2mPipe_rData_twiceMode;
  wire                when_Stream_l368_8;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_valid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_ready;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_frameStart;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_rowEnd;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passMode;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passValid;
  wire       [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceMode;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceValid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainCompare;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterCompare;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDiff;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceCompValid;
  wire       [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceMode;
  reg                 controlStream_s2mPipe_m2sPipe_rValid;
  reg                 controlStream_s2mPipe_m2sPipe_rData_frameStart;
  reg                 controlStream_s2mPipe_m2sPipe_rData_rowEnd;
  reg                 controlStream_s2mPipe_m2sPipe_rData_passMode;
  reg                 controlStream_s2mPipe_m2sPipe_rData_passValid;
  reg        [2:0]    controlStream_s2mPipe_m2sPipe_rData_onceMode;
  reg                 controlStream_s2mPipe_m2sPipe_rData_onceValid;
  reg                 controlStream_s2mPipe_m2sPipe_rData_mainCompare;
  reg                 controlStream_s2mPipe_m2sPipe_rData_counterCompare;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_rData_mainDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_rData_counterDiff;
  reg                 controlStream_s2mPipe_m2sPipe_rData_twiceCompValid;
  reg        [2:0]    controlStream_s2mPipe_m2sPipe_rData_twiceMode;
  wire                when_Stream_l368_9;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_valid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_frameStart;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_rowEnd;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_passMode;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_passValid;
  wire       [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_onceMode;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_onceValid;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainCompare;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterCompare;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainDiff;
  wire       [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterDiff;
  wire                controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_twiceCompValid;
  wire       [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_twiceMode;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_frameStart;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_rowEnd;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_passMode;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_passValid;
  reg        [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_onceMode;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_onceValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainCompare;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterCompare;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterDiff;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_rData_twiceCompValid;
  reg        [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_rData_twiceMode;
  wire                readStage_controlPipe_valid;
  wire                readStage_controlPipe_ready;
  wire                readStage_controlPipe_payload_frameStart;
  wire                readStage_controlPipe_payload_rowEnd;
  wire                readStage_controlPipe_payload_passMode;
  wire                readStage_controlPipe_payload_passValid;
  wire       [2:0]    readStage_controlPipe_payload_onceMode;
  wire                readStage_controlPipe_payload_onceValid;
  wire                readStage_controlPipe_payload_mainCompare;
  wire                readStage_controlPipe_payload_counterCompare;
  wire       [7:0]    readStage_controlPipe_payload_mainDiff;
  wire       [7:0]    readStage_controlPipe_payload_counterDiff;
  wire                readStage_controlPipe_payload_twiceCompValid;
  wire       [2:0]    readStage_controlPipe_payload_twiceMode;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_frameStart;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_rowEnd;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_passMode;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_passValid;
  reg        [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_onceMode;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_onceValid;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainCompare;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterCompare;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainDiff;
  reg        [7:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterDiff;
  reg                 controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_twiceCompValid;
  reg        [2:0]    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_twiceMode;
  wire                when_Stream_l368_10;
  wire                readStage_mainOnePixelStream_s2mPipe_valid;
  reg                 readStage_mainOnePixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_mainOnePixelStream_s2mPipe_payload;
  reg                 readStage_mainOnePixelStream_rValid;
  reg        [7:0]    readStage_mainOnePixelStream_rData;
  wire                compareStage_mainOnePixelStream_valid;
  wire                compareStage_mainOnePixelStream_ready;
  wire       [7:0]    compareStage_mainOnePixelStream_payload;
  reg                 readStage_mainOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_mainOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_11;
  wire                readStage_counterOnePixelStream_s2mPipe_valid;
  reg                 readStage_counterOnePixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_counterOnePixelStream_s2mPipe_payload;
  reg                 readStage_counterOnePixelStream_rValid;
  reg        [7:0]    readStage_counterOnePixelStream_rData;
  wire                compareStage_counterOnePixelStream_valid;
  wire                compareStage_counterOnePixelStream_ready;
  wire       [7:0]    compareStage_counterOnePixelStream_payload;
  reg                 readStage_counterOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_counterOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_12;
  wire                readStage_mainTwoPixelStream_s2mPipe_valid;
  reg                 readStage_mainTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_mainTwoPixelStream_s2mPipe_payload;
  reg                 readStage_mainTwoPixelStream_rValid;
  reg        [7:0]    readStage_mainTwoPixelStream_rData;
  wire                compareStage_mainTwoPixelStream_valid;
  wire                compareStage_mainTwoPixelStream_ready;
  wire       [7:0]    compareStage_mainTwoPixelStream_payload;
  reg                 readStage_mainTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_mainTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_13;
  wire                readStage_counterTwoPixelStream_s2mPipe_valid;
  reg                 readStage_counterTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    readStage_counterTwoPixelStream_s2mPipe_payload;
  reg                 readStage_counterTwoPixelStream_rValid;
  reg        [7:0]    readStage_counterTwoPixelStream_rData;
  wire                compareStage_counterTwoPixelStream_valid;
  wire                compareStage_counterTwoPixelStream_ready;
  wire       [7:0]    compareStage_counterTwoPixelStream_payload;
  reg                 readStage_counterTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    readStage_counterTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_14;
  reg                 CICC1851_readStage_controlPipe_translated_payload_mainCompare;
  reg                 CICC1851_readStage_controlPipe_translated_payload_counterCompare;
  wire                when_SuperResolutionPart1_l205;
  wire                when_SuperResolutionPart1_l209;
  wire                when_SuperResolutionPart1_l213;
  wire                when_SuperResolutionPart1_l217;
  wire                when_SuperResolutionPart1_l228;
  wire                when_SuperResolutionPart1_l230;
  wire                when_SuperResolutionPart1_l234;
  wire                when_SuperResolutionPart1_l236;
  wire                when_SuperResolutionPart1_l241;
  wire                when_SuperResolutionPart1_l246;
  wire                readStage_controlPipe_translated_valid;
  wire                readStage_controlPipe_translated_ready;
  wire                readStage_controlPipe_translated_payload_frameStart;
  wire                readStage_controlPipe_translated_payload_rowEnd;
  wire                readStage_controlPipe_translated_payload_passMode;
  wire                readStage_controlPipe_translated_payload_passValid;
  wire       [2:0]    readStage_controlPipe_translated_payload_onceMode;
  wire                readStage_controlPipe_translated_payload_onceValid;
  wire                readStage_controlPipe_translated_payload_mainCompare;
  wire                readStage_controlPipe_translated_payload_counterCompare;
  wire       [7:0]    readStage_controlPipe_translated_payload_mainDiff;
  wire       [7:0]    readStage_controlPipe_translated_payload_counterDiff;
  wire                readStage_controlPipe_translated_payload_twiceCompValid;
  wire       [2:0]    readStage_controlPipe_translated_payload_twiceMode;
  wire                readStage_controlPipe_translated_s2mPipe_valid;
  reg                 readStage_controlPipe_translated_s2mPipe_ready;
  wire                readStage_controlPipe_translated_s2mPipe_payload_frameStart;
  wire                readStage_controlPipe_translated_s2mPipe_payload_rowEnd;
  wire                readStage_controlPipe_translated_s2mPipe_payload_passMode;
  wire                readStage_controlPipe_translated_s2mPipe_payload_passValid;
  wire       [2:0]    readStage_controlPipe_translated_s2mPipe_payload_onceMode;
  wire                readStage_controlPipe_translated_s2mPipe_payload_onceValid;
  wire                readStage_controlPipe_translated_s2mPipe_payload_mainCompare;
  wire                readStage_controlPipe_translated_s2mPipe_payload_counterCompare;
  wire       [7:0]    readStage_controlPipe_translated_s2mPipe_payload_mainDiff;
  wire       [7:0]    readStage_controlPipe_translated_s2mPipe_payload_counterDiff;
  wire                readStage_controlPipe_translated_s2mPipe_payload_twiceCompValid;
  wire       [2:0]    readStage_controlPipe_translated_s2mPipe_payload_twiceMode;
  reg                 readStage_controlPipe_translated_rValid;
  reg                 readStage_controlPipe_translated_rData_frameStart;
  reg                 readStage_controlPipe_translated_rData_rowEnd;
  reg                 readStage_controlPipe_translated_rData_passMode;
  reg                 readStage_controlPipe_translated_rData_passValid;
  reg        [2:0]    readStage_controlPipe_translated_rData_onceMode;
  reg                 readStage_controlPipe_translated_rData_onceValid;
  reg                 readStage_controlPipe_translated_rData_mainCompare;
  reg                 readStage_controlPipe_translated_rData_counterCompare;
  reg        [7:0]    readStage_controlPipe_translated_rData_mainDiff;
  reg        [7:0]    readStage_controlPipe_translated_rData_counterDiff;
  reg                 readStage_controlPipe_translated_rData_twiceCompValid;
  reg        [2:0]    readStage_controlPipe_translated_rData_twiceMode;
  wire                compareStage_controlPipe_valid;
  wire                compareStage_controlPipe_ready;
  wire                compareStage_controlPipe_payload_frameStart;
  wire                compareStage_controlPipe_payload_rowEnd;
  wire                compareStage_controlPipe_payload_passMode;
  wire                compareStage_controlPipe_payload_passValid;
  wire       [2:0]    compareStage_controlPipe_payload_onceMode;
  wire                compareStage_controlPipe_payload_onceValid;
  wire                compareStage_controlPipe_payload_mainCompare;
  wire                compareStage_controlPipe_payload_counterCompare;
  wire       [7:0]    compareStage_controlPipe_payload_mainDiff;
  wire       [7:0]    compareStage_controlPipe_payload_counterDiff;
  wire                compareStage_controlPipe_payload_twiceCompValid;
  wire       [2:0]    compareStage_controlPipe_payload_twiceMode;
  reg                 readStage_controlPipe_translated_s2mPipe_rValid;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_frameStart;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_rowEnd;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_passMode;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_passValid;
  reg        [2:0]    readStage_controlPipe_translated_s2mPipe_rData_onceMode;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_onceValid;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_mainCompare;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_counterCompare;
  reg        [7:0]    readStage_controlPipe_translated_s2mPipe_rData_mainDiff;
  reg        [7:0]    readStage_controlPipe_translated_s2mPipe_rData_counterDiff;
  reg                 readStage_controlPipe_translated_s2mPipe_rData_twiceCompValid;
  reg        [2:0]    readStage_controlPipe_translated_s2mPipe_rData_twiceMode;
  wire                when_Stream_l368_15;
  wire                compareStage_mainOnePixelStream_s2mPipe_valid;
  reg                 compareStage_mainOnePixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_mainOnePixelStream_s2mPipe_payload;
  reg                 compareStage_mainOnePixelStream_rValid;
  reg        [7:0]    compareStage_mainOnePixelStream_rData;
  wire                diffStage_mainOnePixelStream_valid;
  wire                diffStage_mainOnePixelStream_ready;
  wire       [7:0]    diffStage_mainOnePixelStream_payload;
  reg                 compareStage_mainOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_mainOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_16;
  wire                compareStage_counterOnePixelStream_s2mPipe_valid;
  reg                 compareStage_counterOnePixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_counterOnePixelStream_s2mPipe_payload;
  reg                 compareStage_counterOnePixelStream_rValid;
  reg        [7:0]    compareStage_counterOnePixelStream_rData;
  wire                diffStage_counterOnePixelStream_valid;
  wire                diffStage_counterOnePixelStream_ready;
  wire       [7:0]    diffStage_counterOnePixelStream_payload;
  reg                 compareStage_counterOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_counterOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_17;
  wire                compareStage_mainTwoPixelStream_s2mPipe_valid;
  reg                 compareStage_mainTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_mainTwoPixelStream_s2mPipe_payload;
  reg                 compareStage_mainTwoPixelStream_rValid;
  reg        [7:0]    compareStage_mainTwoPixelStream_rData;
  wire                diffStage_mainTwoPixelStream_valid;
  wire                diffStage_mainTwoPixelStream_ready;
  wire       [7:0]    diffStage_mainTwoPixelStream_payload;
  reg                 compareStage_mainTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_mainTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_18;
  wire                compareStage_counterTwoPixelStream_s2mPipe_valid;
  reg                 compareStage_counterTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    compareStage_counterTwoPixelStream_s2mPipe_payload;
  reg                 compareStage_counterTwoPixelStream_rValid;
  reg        [7:0]    compareStage_counterTwoPixelStream_rData;
  wire                diffStage_counterTwoPixelStream_valid;
  wire                diffStage_counterTwoPixelStream_ready;
  wire       [7:0]    diffStage_counterTwoPixelStream_payload;
  reg                 compareStage_counterTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    compareStage_counterTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_19;
  reg        [7:0]    CICC1851_compareStage_controlPipe_translated_payload_mainDiff;
  reg        [7:0]    CICC1851_compareStage_controlPipe_translated_payload_counterDiff;
  wire                compareStage_controlPipe_translated_valid;
  wire                compareStage_controlPipe_translated_ready;
  wire                compareStage_controlPipe_translated_payload_frameStart;
  wire                compareStage_controlPipe_translated_payload_rowEnd;
  wire                compareStage_controlPipe_translated_payload_passMode;
  wire                compareStage_controlPipe_translated_payload_passValid;
  wire       [2:0]    compareStage_controlPipe_translated_payload_onceMode;
  wire                compareStage_controlPipe_translated_payload_onceValid;
  wire                compareStage_controlPipe_translated_payload_mainCompare;
  wire                compareStage_controlPipe_translated_payload_counterCompare;
  wire       [7:0]    compareStage_controlPipe_translated_payload_mainDiff;
  wire       [7:0]    compareStage_controlPipe_translated_payload_counterDiff;
  wire                compareStage_controlPipe_translated_payload_twiceCompValid;
  wire       [2:0]    compareStage_controlPipe_translated_payload_twiceMode;
  wire                compareStage_controlPipe_translated_s2mPipe_valid;
  reg                 compareStage_controlPipe_translated_s2mPipe_ready;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_frameStart;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_rowEnd;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_passMode;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_passValid;
  wire       [2:0]    compareStage_controlPipe_translated_s2mPipe_payload_onceMode;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_onceValid;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_mainCompare;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_counterCompare;
  wire       [7:0]    compareStage_controlPipe_translated_s2mPipe_payload_mainDiff;
  wire       [7:0]    compareStage_controlPipe_translated_s2mPipe_payload_counterDiff;
  wire                compareStage_controlPipe_translated_s2mPipe_payload_twiceCompValid;
  wire       [2:0]    compareStage_controlPipe_translated_s2mPipe_payload_twiceMode;
  reg                 compareStage_controlPipe_translated_rValid;
  reg                 compareStage_controlPipe_translated_rData_frameStart;
  reg                 compareStage_controlPipe_translated_rData_rowEnd;
  reg                 compareStage_controlPipe_translated_rData_passMode;
  reg                 compareStage_controlPipe_translated_rData_passValid;
  reg        [2:0]    compareStage_controlPipe_translated_rData_onceMode;
  reg                 compareStage_controlPipe_translated_rData_onceValid;
  reg                 compareStage_controlPipe_translated_rData_mainCompare;
  reg                 compareStage_controlPipe_translated_rData_counterCompare;
  reg        [7:0]    compareStage_controlPipe_translated_rData_mainDiff;
  reg        [7:0]    compareStage_controlPipe_translated_rData_counterDiff;
  reg                 compareStage_controlPipe_translated_rData_twiceCompValid;
  reg        [2:0]    compareStage_controlPipe_translated_rData_twiceMode;
  wire                diffStage_controlPipe_valid;
  wire                diffStage_controlPipe_ready;
  wire                diffStage_controlPipe_payload_frameStart;
  wire                diffStage_controlPipe_payload_rowEnd;
  wire                diffStage_controlPipe_payload_passMode;
  wire                diffStage_controlPipe_payload_passValid;
  wire       [2:0]    diffStage_controlPipe_payload_onceMode;
  wire                diffStage_controlPipe_payload_onceValid;
  wire                diffStage_controlPipe_payload_mainCompare;
  wire                diffStage_controlPipe_payload_counterCompare;
  wire       [7:0]    diffStage_controlPipe_payload_mainDiff;
  wire       [7:0]    diffStage_controlPipe_payload_counterDiff;
  wire                diffStage_controlPipe_payload_twiceCompValid;
  wire       [2:0]    diffStage_controlPipe_payload_twiceMode;
  reg                 compareStage_controlPipe_translated_s2mPipe_rValid;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_frameStart;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_rowEnd;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_passMode;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_passValid;
  reg        [2:0]    compareStage_controlPipe_translated_s2mPipe_rData_onceMode;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_onceValid;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_mainCompare;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_counterCompare;
  reg        [7:0]    compareStage_controlPipe_translated_s2mPipe_rData_mainDiff;
  reg        [7:0]    compareStage_controlPipe_translated_s2mPipe_rData_counterDiff;
  reg                 compareStage_controlPipe_translated_s2mPipe_rData_twiceCompValid;
  reg        [2:0]    compareStage_controlPipe_translated_s2mPipe_rData_twiceMode;
  wire                when_Stream_l368_20;
  wire                diffStage_mainOnePixelStream_s2mPipe_valid;
  reg                 diffStage_mainOnePixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_mainOnePixelStream_s2mPipe_payload;
  reg                 diffStage_mainOnePixelStream_rValid;
  reg        [7:0]    diffStage_mainOnePixelStream_rData;
  wire                resultStage_mainOnePixelStream_valid;
  wire                resultStage_mainOnePixelStream_ready;
  wire       [7:0]    resultStage_mainOnePixelStream_payload;
  reg                 diffStage_mainOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_mainOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_21;
  wire                diffStage_counterOnePixelStream_s2mPipe_valid;
  reg                 diffStage_counterOnePixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_counterOnePixelStream_s2mPipe_payload;
  reg                 diffStage_counterOnePixelStream_rValid;
  reg        [7:0]    diffStage_counterOnePixelStream_rData;
  wire                resultStage_counterOnePixelStream_valid;
  wire                resultStage_counterOnePixelStream_ready;
  wire       [7:0]    resultStage_counterOnePixelStream_payload;
  reg                 diffStage_counterOnePixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_counterOnePixelStream_s2mPipe_rData;
  wire                when_Stream_l368_22;
  wire                diffStage_mainTwoPixelStream_s2mPipe_valid;
  reg                 diffStage_mainTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_mainTwoPixelStream_s2mPipe_payload;
  reg                 diffStage_mainTwoPixelStream_rValid;
  reg        [7:0]    diffStage_mainTwoPixelStream_rData;
  wire                resultStage_mainTwoPixelStream_valid;
  wire                resultStage_mainTwoPixelStream_ready;
  wire       [7:0]    resultStage_mainTwoPixelStream_payload;
  reg                 diffStage_mainTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_mainTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_23;
  wire                diffStage_counterTwoPixelStream_s2mPipe_valid;
  reg                 diffStage_counterTwoPixelStream_s2mPipe_ready;
  wire       [7:0]    diffStage_counterTwoPixelStream_s2mPipe_payload;
  reg                 diffStage_counterTwoPixelStream_rValid;
  reg        [7:0]    diffStage_counterTwoPixelStream_rData;
  wire                resultStage_counterTwoPixelStream_valid;
  wire                resultStage_counterTwoPixelStream_ready;
  wire       [7:0]    resultStage_counterTwoPixelStream_payload;
  reg                 diffStage_counterTwoPixelStream_s2mPipe_rValid;
  reg        [7:0]    diffStage_counterTwoPixelStream_s2mPipe_rData;
  wire                when_Stream_l368_24;
  wire                diffStage_controlPipe_fork_io_outputs_0_s2mPipe_valid;
  reg                 diffStage_controlPipe_fork_io_outputs_0_s2mPipe_ready;
  wire                diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_frameStart;
  wire                diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_rowEnd;
  wire                diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_passMode;
  wire                diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_passValid;
  wire       [2:0]    diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_onceMode;
  wire                diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_onceValid;
  wire                diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_mainCompare;
  wire                diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_counterCompare;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_mainDiff;
  wire       [7:0]    diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_counterDiff;
  wire                diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_twiceCompValid;
  wire       [2:0]    diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_twiceMode;
  reg                 diffStage_controlPipe_fork_io_outputs_0_rValid;
  reg                 diffStage_controlPipe_fork_io_outputs_0_rData_frameStart;
  reg                 diffStage_controlPipe_fork_io_outputs_0_rData_rowEnd;
  reg                 diffStage_controlPipe_fork_io_outputs_0_rData_passMode;
  reg                 diffStage_controlPipe_fork_io_outputs_0_rData_passValid;
  reg        [2:0]    diffStage_controlPipe_fork_io_outputs_0_rData_onceMode;
  reg                 diffStage_controlPipe_fork_io_outputs_0_rData_onceValid;
  reg                 diffStage_controlPipe_fork_io_outputs_0_rData_mainCompare;
  reg                 diffStage_controlPipe_fork_io_outputs_0_rData_counterCompare;
  reg        [7:0]    diffStage_controlPipe_fork_io_outputs_0_rData_mainDiff;
  reg        [7:0]    diffStage_controlPipe_fork_io_outputs_0_rData_counterDiff;
  reg                 diffStage_controlPipe_fork_io_outputs_0_rData_twiceCompValid;
  reg        [2:0]    diffStage_controlPipe_fork_io_outputs_0_rData_twiceMode;
  wire                resultStage_controlPipe_valid;
  wire                resultStage_controlPipe_ready;
  wire                resultStage_controlPipe_payload_frameStart;
  wire                resultStage_controlPipe_payload_rowEnd;
  wire                resultStage_controlPipe_payload_passMode;
  wire                resultStage_controlPipe_payload_passValid;
  wire       [2:0]    resultStage_controlPipe_payload_onceMode;
  wire                resultStage_controlPipe_payload_onceValid;
  wire                resultStage_controlPipe_payload_mainCompare;
  wire                resultStage_controlPipe_payload_counterCompare;
  wire       [7:0]    resultStage_controlPipe_payload_mainDiff;
  wire       [7:0]    resultStage_controlPipe_payload_counterDiff;
  wire                resultStage_controlPipe_payload_twiceCompValid;
  wire       [2:0]    resultStage_controlPipe_payload_twiceMode;
  reg                 diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rValid;
  reg                 diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_frameStart;
  reg                 diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_rowEnd;
  reg                 diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_passMode;
  reg                 diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_passValid;
  reg        [2:0]    diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_onceMode;
  reg                 diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_onceValid;
  reg                 diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_mainCompare;
  reg                 diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_counterCompare;
  reg        [7:0]    diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_mainDiff;
  reg        [7:0]    diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_counterDiff;
  reg                 diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_twiceCompValid;
  reg        [2:0]    diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_twiceMode;
  wire                when_Stream_l368_25;
  wire                resultStage_pixelStream_valid;
  wire                resultStage_pixelStream_ready;
  reg        [7:0]    resultStage_pixelStream_payload;
  wire                when_SuperResolutionPart1_l339;
  wire                when_SuperResolutionPart1_l343;
  wire                when_SuperResolutionPart1_l347;
  wire                when_SuperResolutionPart1_l351;
  wire                when_SuperResolutionPart1_l362;
  wire                when_SuperResolutionPart1_l363;
  wire                when_SuperResolutionPart1_l366;
  wire                when_SuperResolutionPart1_l371;
  wire                when_SuperResolutionPart1_l372;
  wire                when_SuperResolutionPart1_l375;
  wire                when_SuperResolutionPart1_l381;
  wire                when_SuperResolutionPart1_l386;
  wire                resultStage_pixelStream_s2mPipe_valid;
  reg                 resultStage_pixelStream_s2mPipe_ready;
  wire       [7:0]    resultStage_pixelStream_s2mPipe_payload;
  reg                 resultStage_pixelStream_rValid;
  reg        [7:0]    resultStage_pixelStream_rData;
  wire                resultStage_resultStream_valid;
  wire                resultStage_resultStream_ready;
  wire       [7:0]    resultStage_resultStream_payload;
  reg                 resultStage_pixelStream_s2mPipe_rValid;
  reg        [7:0]    resultStage_pixelStream_s2mPipe_rData;
  wire                when_Stream_l368_26;
  wire                CICC1851_resultStage_mainOnePixelStream_ready;
  reg                 CICC1851_resultStage_mainOnePixelStream_ready_1;
  wire                CICC1851_resultStage_mainOnePixelStream_ready_2;
  wire                when_Stream_l438;
  reg                 resultsJoin_valid;
  wire                resultsJoin_ready;
  wire                pixelsStream_valid;
  wire                pixelsStream_ready;
  wire       [7:0]    pixelsStream_payload_pixel;
  wire                pixelsStream_payload_frameStart;
  wire                pixelsStream_payload_rowEnd;
  wire                pixelsStream_s2mPipe_valid;
  reg                 pixelsStream_s2mPipe_ready;
  wire       [7:0]    pixelsStream_s2mPipe_payload_pixel;
  wire                pixelsStream_s2mPipe_payload_frameStart;
  wire                pixelsStream_s2mPipe_payload_rowEnd;
  reg                 pixelsStream_rValid;
  reg        [7:0]    pixelsStream_rData_pixel;
  reg                 pixelsStream_rData_frameStart;
  reg                 pixelsStream_rData_rowEnd;
  wire                pixelsStream_s2mPipe_m2sPipe_valid;
  wire                pixelsStream_s2mPipe_m2sPipe_ready;
  wire       [7:0]    pixelsStream_s2mPipe_m2sPipe_payload_pixel;
  wire                pixelsStream_s2mPipe_m2sPipe_payload_frameStart;
  wire                pixelsStream_s2mPipe_m2sPipe_payload_rowEnd;
  reg                 pixelsStream_s2mPipe_rValid;
  reg        [7:0]    pixelsStream_s2mPipe_rData_pixel;
  reg                 pixelsStream_s2mPipe_rData_frameStart;
  reg                 pixelsStream_s2mPipe_rData_rowEnd;
  wire                when_Stream_l368_27;
  wire                pixelsIn_s2mPipe_valid;
  reg                 pixelsIn_s2mPipe_ready;
  wire       [7:0]    pixelsIn_s2mPipe_payload_pixel;
  wire                pixelsIn_s2mPipe_payload_frameStart;
  wire                pixelsIn_s2mPipe_payload_rowEnd;
  reg                 pixelsIn_rValid;
  reg        [7:0]    pixelsIn_rData_pixel;
  reg                 pixelsIn_rData_frameStart;
  reg                 pixelsIn_rData_rowEnd;
  wire                pixelsIn_s2mPipe_m2sPipe_valid;
  wire                pixelsIn_s2mPipe_m2sPipe_ready;
  wire       [7:0]    pixelsIn_s2mPipe_m2sPipe_payload_pixel;
  wire                pixelsIn_s2mPipe_m2sPipe_payload_frameStart;
  wire                pixelsIn_s2mPipe_m2sPipe_payload_rowEnd;
  reg                 pixelsIn_s2mPipe_rValid;
  reg        [7:0]    pixelsIn_s2mPipe_rData_pixel;
  reg                 pixelsIn_s2mPipe_rData_frameStart;
  reg                 pixelsIn_s2mPipe_rData_rowEnd;
  wire                when_Stream_l368_28;
  wire                passPixels_valid;
  wire                passPixels_ready;
  wire       [7:0]    passPixels_payload_pixel;
  wire                passPixels_payload_frameStart;
  wire                passPixels_payload_rowEnd;
  wire                passPixels_fire;
  wire                when_SuperResolutionPart1_l421;
  wire                passPixels_fire_1;
  wire                when_SuperResolutionPart1_l422;
  wire                passPixels_fire_2;
  wire                when_SuperResolutionPart1_l425;
  wire                passPixels_fire_3;
  wire                when_SuperResolutionPart1_l438;
  wire                passPixels_fire_4;
  wire                when_SuperResolutionPart1_l439;
  wire                when_SuperResolutionPart1_l442;
  wire                controlStream_fire;
  wire                when_SuperResolutionPart1_l447;
  wire                when_SuperResolutionPart1_l449;
  wire                passPixels_fire_5;
  wire                when_SuperResolutionPart1_l453;
  wire                passPixels_fire_6;
  wire                passPixels_fire_7;
  wire                passPixels_fire_8;
  wire                controlStateMachine_wantExit;
  reg                 controlStateMachine_wantStart;
  wire                controlStateMachine_wantKill;
  reg        [2:0]    controlStateMachine_stateReg;
  reg        [2:0]    controlStateMachine_stateNext;
  wire                when_SuperResolutionPart1_l482;
  wire                passPixels_fire_9;
  wire                when_SuperResolutionPart1_l484;
  wire                passPixels_fire_10;
  wire                when_SuperResolutionPart1_l489;
  wire                controlStream_fire_1;
  wire                when_SuperResolutionPart1_l498;
  wire                passPixels_fire_11;
  wire                when_SuperResolutionPart1_l500;
  wire                controlStream_fire_2;
  wire                when_SuperResolutionPart1_l507;
  wire                controlStream_fire_3;
  wire                when_SuperResolutionPart1_l510;
  wire                controlStream_fire_4;
  wire                when_SuperResolutionPart1_l511;
  wire                controlStream_fire_5;
  wire                when_SuperResolutionPart1_l513;
  wire                controlStream_fire_6;
  wire                when_SuperResolutionPart1_l537;
  wire                controlStream_fire_7;
  wire                when_SuperResolutionPart1_l542;
  wire                controlStream_fire_8;
  wire                passPixels_fire_12;
  wire                when_SuperResolutionPart1_l563;
  wire                controlStream_fire_9;
  wire                when_SuperResolutionPart1_l578;
  wire                controlStream_fire_10;
  wire                when_SuperResolutionPart1_l579;
  wire                controlStream_fire_11;
  wire                when_SuperResolutionPart1_l581;
  wire                controlStream_fire_12;
  wire                controlStream_fire_13;
  wire                when_SuperResolutionPart1_l612;
  wire                controlStream_fire_14;
  wire                when_SuperResolutionPart1_l664;
  wire                controlStream_fire_15;
  wire                when_SuperResolutionPart1_l665;
  wire                controlStream_fire_16;
  wire                when_SuperResolutionPart1_l667;
  wire                controlStream_fire_17;
  `ifndef SYNTHESIS
  reg [39:0] controlStateMachine_stateReg_string;
  reg [39:0] controlStateMachine_stateNext_string;
  `endif

  reg [7:0] lineBufferOne [0:959];
  reg [7:0] lineBufferTwo [0:959];

  assign CICC1851_bufferRowCount_valueNext_1 = bufferRowCount_willIncrement;
  assign CICC1851_bufferRowCount_valueNext = {9'd0, CICC1851_bufferRowCount_valueNext_1};
  assign CICC1851_bufferWAddr_valueNext_1 = bufferWAddr_willIncrement;
  assign CICC1851_bufferWAddr_valueNext = {9'd0, CICC1851_bufferWAddr_valueNext_1};
  assign CICC1851_outPixelAddr_valueNext_1 = outPixelAddr_willIncrement;
  assign CICC1851_outPixelAddr_valueNext = {10'd0, CICC1851_outPixelAddr_valueNext_1};
  assign CICC1851_outRowCount_valueNext_1 = outRowCount_willIncrement;
  assign CICC1851_outRowCount_valueNext = {10'd0, CICC1851_outRowCount_valueNext_1};
  assign CICC1851_mainAddrOne = (outPixelAddr_value / 2'b10);
  assign CICC1851_counterAddrOne = (outPixelAddr_value / 2'b10);
  assign CICC1851_mainAddrTwo = (outPixelAddr_value / 2'b10);
  assign CICC1851_counterAddrTwo = (outPixelAddr_value / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload = (CICC1851_resultStage_pixelStream_payload_1 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_1 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_2 = (CICC1851_resultStage_pixelStream_payload_3 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_3 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_4 = (CICC1851_resultStage_pixelStream_payload_5 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_5 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_mainTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_6 = (CICC1851_resultStage_pixelStream_payload_7 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_7 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_mainOnePixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_8 = (CICC1851_resultStage_pixelStream_payload_9 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_9 = ({1'b0,diffStage_counterOnePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_10 = (CICC1851_resultStage_pixelStream_payload_11 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_11 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_mainTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_12 = (CICC1851_resultStage_pixelStream_payload_13 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_13 = ({1'b0,diffStage_counterOnePixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_14 = (CICC1851_resultStage_pixelStream_payload_15 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_15 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_mainTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_16 = (CICC1851_resultStage_pixelStream_payload_17 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_17 = ({1'b0,diffStage_mainTwoPixelStream_payload} + {1'b0,diffStage_counterTwoPixelStream_payload});
  assign CICC1851_resultStage_pixelStream_payload_18 = (CICC1851_resultStage_pixelStream_payload_19 / 2'b10);
  assign CICC1851_resultStage_pixelStream_payload_19 = ({1'b0,diffStage_mainOnePixelStream_payload} + {1'b0,diffStage_counterOnePixelStream_payload});
  assign CICC1851_when_SuperResolutionPart1_l421 = (bmpWidth - 10'h002);
  assign CICC1851_when_SuperResolutionPart1_l422 = (bmpHeight - 10'h002);
  assign CICC1851_when_SuperResolutionPart1_l447 = (outRowCount_value % 2'b10);
  assign CICC1851_when_SuperResolutionPart1_l482 = (outRowCount_value % 2'b10);
  assign CICC1851_when_SuperResolutionPart1_l484 = (outPixelAddr_value % 2'b10);
  assign CICC1851_when_SuperResolutionPart1_l489 = (outPixelAddr_value % 2'b10);
  assign CICC1851_when_SuperResolutionPart1_l498 = {1'd0, outRowCount_value};
  assign CICC1851_when_SuperResolutionPart1_l498_1 = (2'b10 * bufferRowCount_value);
  assign CICC1851_when_SuperResolutionPart1_l500 = (2'b10 * bufferWAddr_value);
  assign CICC1851_when_SuperResolutionPart1_l500_1 = ({1'b0,outPixelAddr_value} + CICC1851_when_SuperResolutionPart1_l500_2);
  assign CICC1851_when_SuperResolutionPart1_l500_3 = {1'b0,2'b10};
  assign CICC1851_when_SuperResolutionPart1_l500_2 = {9'd0, CICC1851_when_SuperResolutionPart1_l500_3};
  assign CICC1851_when_SuperResolutionPart1_l510 = {1'd0, outPixelAddr_value};
  assign CICC1851_when_SuperResolutionPart1_l510_1 = (CICC1851_when_SuperResolutionPart1_l510_2 - 12'h002);
  assign CICC1851_when_SuperResolutionPart1_l510_2 = (2'b10 * bmpWidth);
  assign CICC1851_when_SuperResolutionPart1_l511 = {1'd0, outRowCount_value};
  assign CICC1851_when_SuperResolutionPart1_l511_1 = (CICC1851_when_SuperResolutionPart1_l511_2 - 12'h002);
  assign CICC1851_when_SuperResolutionPart1_l511_2 = (2'b10 * bmpHeight);
  assign CICC1851_when_SuperResolutionPart1_l537 = (outRowCount_value % 2'b10);
  assign CICC1851_when_SuperResolutionPart1_l542_1 = (11'h002 + outRowCount_value);
  assign CICC1851_when_SuperResolutionPart1_l542 = {1'd0, CICC1851_when_SuperResolutionPart1_l542_1};
  assign CICC1851_when_SuperResolutionPart1_l542_2 = (2'b10 * bufferRowCount_value);
  assign CICC1851_mainAddrOne_1 = (CICC1851_mainAddrOne_2 / 2'b10);
  assign CICC1851_mainAddrOne_2 = (outPixelAddr_value - 11'h001);
  assign CICC1851_counterAddrOne_1 = (CICC1851_counterAddrOne_2 / 2'b10);
  assign CICC1851_counterAddrOne_2 = (outPixelAddr_value - 11'h001);
  assign CICC1851_counterAddrOne_3 = (CICC1851_counterAddrOne_4 / 2'b10);
  assign CICC1851_counterAddrOne_4 = ({1'b0,outPixelAddr_value} + CICC1851_counterAddrOne_5);
  assign CICC1851_counterAddrOne_6 = {1'b0,1'b1};
  assign CICC1851_counterAddrOne_5 = {10'd0, CICC1851_counterAddrOne_6};
  assign CICC1851_controls_onceMode = 1'b1;
  assign CICC1851_mainAddrTwo_1 = (CICC1851_mainAddrTwo_2 / 2'b10);
  assign CICC1851_mainAddrTwo_2 = (outPixelAddr_value - 11'h001);
  assign CICC1851_counterAddrTwo_1 = (CICC1851_counterAddrTwo_2 / 2'b10);
  assign CICC1851_counterAddrTwo_2 = (outPixelAddr_value - 11'h001);
  assign CICC1851_counterAddrTwo_3 = (CICC1851_counterAddrTwo_4 / 2'b10);
  assign CICC1851_counterAddrTwo_4 = ({1'b0,outPixelAddr_value} + CICC1851_counterAddrTwo_5);
  assign CICC1851_counterAddrTwo_6 = {1'b0,1'b1};
  assign CICC1851_counterAddrTwo_5 = {10'd0, CICC1851_counterAddrTwo_6};
  assign CICC1851_when_SuperResolutionPart1_l563 = (2'b10 * bufferWAddr_value);
  assign CICC1851_when_SuperResolutionPart1_l563_1 = ({1'b0,outPixelAddr_value} + CICC1851_when_SuperResolutionPart1_l563_2);
  assign CICC1851_when_SuperResolutionPart1_l563_3 = {1'b0,2'b10};
  assign CICC1851_when_SuperResolutionPart1_l563_2 = {9'd0, CICC1851_when_SuperResolutionPart1_l563_3};
  assign CICC1851_controls_onceMode_1 = 2'b10;
  assign CICC1851_controls_onceMode_2 = 2'b11;
  assign CICC1851_mainAddrOne_3 = (outPixelAddr_value / 2'b10);
  assign CICC1851_mainAddrTwo_3 = (outPixelAddr_value / 2'b10);
  assign CICC1851_when_SuperResolutionPart1_l578 = {1'd0, outPixelAddr_value};
  assign CICC1851_when_SuperResolutionPart1_l578_1 = (CICC1851_when_SuperResolutionPart1_l578_2 - 12'h002);
  assign CICC1851_when_SuperResolutionPart1_l578_2 = (2'b10 * bmpWidth);
  assign CICC1851_when_SuperResolutionPart1_l579 = {1'd0, outRowCount_value};
  assign CICC1851_when_SuperResolutionPart1_l579_1 = (CICC1851_when_SuperResolutionPart1_l579_2 - 12'h002);
  assign CICC1851_when_SuperResolutionPart1_l579_2 = (2'b10 * bmpHeight);
  assign CICC1851_mainAddrOne_4 = (CICC1851_mainAddrOne_5 / 2'b10);
  assign CICC1851_mainAddrOne_5 = (outPixelAddr_value - 11'h001);
  assign CICC1851_mainAddrOne_6 = (CICC1851_mainAddrOne_7 / 2'b10);
  assign CICC1851_mainAddrOne_7 = (outPixelAddr_value - 11'h001);
  assign CICC1851_counterAddrOne_7 = (CICC1851_counterAddrOne_8 / 2'b10);
  assign CICC1851_counterAddrOne_8 = ({1'b0,outPixelAddr_value} + CICC1851_counterAddrOne_9);
  assign CICC1851_counterAddrOne_10 = {1'b0,1'b1};
  assign CICC1851_counterAddrOne_9 = {10'd0, CICC1851_counterAddrOne_10};
  assign CICC1851_mainAddrTwo_4 = (CICC1851_mainAddrTwo_5 / 2'b10);
  assign CICC1851_mainAddrTwo_5 = (outPixelAddr_value - 11'h001);
  assign CICC1851_mainAddrTwo_6 = (CICC1851_mainAddrTwo_7 / 2'b10);
  assign CICC1851_mainAddrTwo_7 = (outPixelAddr_value - 11'h001);
  assign CICC1851_counterAddrTwo_7 = (CICC1851_counterAddrTwo_8 / 2'b10);
  assign CICC1851_counterAddrTwo_8 = ({1'b0,outPixelAddr_value} + CICC1851_counterAddrTwo_9);
  assign CICC1851_counterAddrTwo_10 = {1'b0,1'b1};
  assign CICC1851_counterAddrTwo_9 = {10'd0, CICC1851_counterAddrTwo_10};
  assign CICC1851_mainAddrOne_8 = (CICC1851_mainAddrOne_9 / 2'b10);
  assign CICC1851_mainAddrOne_9 = (outPixelAddr_value - 11'h001);
  assign CICC1851_counterAddrTwo_11 = (CICC1851_counterAddrTwo_12 / 2'b10);
  assign CICC1851_counterAddrTwo_12 = (outPixelAddr_value - 11'h001);
  assign CICC1851_mainAddrTwo_8 = (CICC1851_mainAddrTwo_9 / 2'b10);
  assign CICC1851_mainAddrTwo_9 = (outPixelAddr_value - 11'h001);
  assign CICC1851_counterAddrOne_11 = (CICC1851_counterAddrOne_12 / 2'b10);
  assign CICC1851_counterAddrOne_12 = (outPixelAddr_value - 11'h001);
  assign CICC1851_mainAddrTwo_10 = (CICC1851_mainAddrTwo_11 / 2'b10);
  assign CICC1851_mainAddrTwo_11 = ({1'b0,outPixelAddr_value} + CICC1851_mainAddrTwo_12);
  assign CICC1851_mainAddrTwo_13 = {1'b0,1'b1};
  assign CICC1851_mainAddrTwo_12 = {10'd0, CICC1851_mainAddrTwo_13};
  assign CICC1851_counterAddrOne_13 = (CICC1851_counterAddrOne_14 / 2'b10);
  assign CICC1851_counterAddrOne_14 = ({1'b0,outPixelAddr_value} + CICC1851_counterAddrOne_15);
  assign CICC1851_counterAddrOne_16 = {1'b0,1'b1};
  assign CICC1851_counterAddrOne_15 = {10'd0, CICC1851_counterAddrOne_16};
  assign CICC1851_mainAddrTwo_14 = (CICC1851_mainAddrTwo_15 / 2'b10);
  assign CICC1851_mainAddrTwo_15 = (outPixelAddr_value - 11'h001);
  assign CICC1851_counterAddrOne_17 = (CICC1851_counterAddrOne_18 / 2'b10);
  assign CICC1851_counterAddrOne_18 = (outPixelAddr_value - 11'h001);
  assign CICC1851_mainAddrOne_10 = (CICC1851_mainAddrOne_11 / 2'b10);
  assign CICC1851_mainAddrOne_11 = (outPixelAddr_value - 11'h001);
  assign CICC1851_counterAddrTwo_13 = (CICC1851_counterAddrTwo_14 / 2'b10);
  assign CICC1851_counterAddrTwo_14 = (outPixelAddr_value - 11'h001);
  assign CICC1851_mainAddrOne_12 = (CICC1851_mainAddrOne_13 / 2'b10);
  assign CICC1851_mainAddrOne_13 = ({1'b0,outPixelAddr_value} + CICC1851_mainAddrOne_14);
  assign CICC1851_mainAddrOne_15 = {1'b0,1'b1};
  assign CICC1851_mainAddrOne_14 = {10'd0, CICC1851_mainAddrOne_15};
  assign CICC1851_counterAddrTwo_15 = (CICC1851_counterAddrTwo_16 / 2'b10);
  assign CICC1851_counterAddrTwo_16 = ({1'b0,outPixelAddr_value} + CICC1851_counterAddrTwo_17);
  assign CICC1851_counterAddrTwo_18 = {1'b0,1'b1};
  assign CICC1851_counterAddrTwo_17 = {10'd0, CICC1851_counterAddrTwo_18};
  assign CICC1851_when_SuperResolutionPart1_l664 = {1'd0, outPixelAddr_value};
  assign CICC1851_when_SuperResolutionPart1_l664_1 = (CICC1851_when_SuperResolutionPart1_l664_2 - 12'h002);
  assign CICC1851_when_SuperResolutionPart1_l664_2 = (2'b10 * bmpWidth);
  assign CICC1851_when_SuperResolutionPart1_l665 = {1'd0, outRowCount_value};
  assign CICC1851_when_SuperResolutionPart1_l665_1 = (CICC1851_when_SuperResolutionPart1_l665_2 - 12'h002);
  assign CICC1851_when_SuperResolutionPart1_l665_2 = (2'b10 * bmpHeight);
  assign CICC1851_lineBufferOne_port = passPixels_payload_pixel;
  assign CICC1851_lineBufferOne_port_1 = (passPixels_fire_7 && (! bufferSwitch));
  assign CICC1851_lineBufferTwo_port = passPixels_payload_pixel;
  assign CICC1851_lineBufferTwo_port_1 = (passPixels_fire_6 && bufferSwitch);
  always @(posedge clk) begin
    if(mainAddrOneStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferOne_port0 <= lineBufferOne[mainAddrOneStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(counterAddrOneStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferOne_port1 <= lineBufferOne[counterAddrOneStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(CICC1851_lineBufferOne_port_1) begin
      lineBufferOne[bufferWAddr_value] <= CICC1851_lineBufferOne_port;
    end
  end

  always @(posedge clk) begin
    if(mainAddrTwoStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferTwo_port0 <= lineBufferTwo[mainAddrTwoStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(counterAddrTwoStream_s2mPipe_m2sPipe_ready) begin
      CICC1851_lineBufferTwo_port1 <= lineBufferTwo[counterAddrTwoStream_s2mPipe_m2sPipe_payload];
    end
  end

  always @(posedge clk) begin
    if(CICC1851_lineBufferTwo_port_1) begin
      lineBufferTwo[bufferWAddr_value] <= CICC1851_lineBufferTwo_port;
    end
  end

  StreamFork_1 diffStage_controlPipe_fork (
    .io_input_valid                      (diffStage_controlPipe_valid                                     ), //i
    .io_input_ready                      (diffStage_controlPipe_fork_io_input_ready                       ), //o
    .io_input_payload_frameStart         (diffStage_controlPipe_payload_frameStart                        ), //i
    .io_input_payload_rowEnd             (diffStage_controlPipe_payload_rowEnd                            ), //i
    .io_input_payload_passMode           (diffStage_controlPipe_payload_passMode                          ), //i
    .io_input_payload_passValid          (diffStage_controlPipe_payload_passValid                         ), //i
    .io_input_payload_onceMode           (diffStage_controlPipe_payload_onceMode[2:0]                     ), //i
    .io_input_payload_onceValid          (diffStage_controlPipe_payload_onceValid                         ), //i
    .io_input_payload_mainCompare        (diffStage_controlPipe_payload_mainCompare                       ), //i
    .io_input_payload_counterCompare     (diffStage_controlPipe_payload_counterCompare                    ), //i
    .io_input_payload_mainDiff           (diffStage_controlPipe_payload_mainDiff[7:0]                     ), //i
    .io_input_payload_counterDiff        (diffStage_controlPipe_payload_counterDiff[7:0]                  ), //i
    .io_input_payload_twiceCompValid     (diffStage_controlPipe_payload_twiceCompValid                    ), //i
    .io_input_payload_twiceMode          (diffStage_controlPipe_payload_twiceMode[2:0]                    ), //i
    .io_outputs_0_valid                  (diffStage_controlPipe_fork_io_outputs_0_valid                   ), //o
    .io_outputs_0_ready                  (diffStage_controlPipe_fork_io_outputs_0_ready                   ), //i
    .io_outputs_0_payload_frameStart     (diffStage_controlPipe_fork_io_outputs_0_payload_frameStart      ), //o
    .io_outputs_0_payload_rowEnd         (diffStage_controlPipe_fork_io_outputs_0_payload_rowEnd          ), //o
    .io_outputs_0_payload_passMode       (diffStage_controlPipe_fork_io_outputs_0_payload_passMode        ), //o
    .io_outputs_0_payload_passValid      (diffStage_controlPipe_fork_io_outputs_0_payload_passValid       ), //o
    .io_outputs_0_payload_onceMode       (diffStage_controlPipe_fork_io_outputs_0_payload_onceMode[2:0]   ), //o
    .io_outputs_0_payload_onceValid      (diffStage_controlPipe_fork_io_outputs_0_payload_onceValid       ), //o
    .io_outputs_0_payload_mainCompare    (diffStage_controlPipe_fork_io_outputs_0_payload_mainCompare     ), //o
    .io_outputs_0_payload_counterCompare (diffStage_controlPipe_fork_io_outputs_0_payload_counterCompare  ), //o
    .io_outputs_0_payload_mainDiff       (diffStage_controlPipe_fork_io_outputs_0_payload_mainDiff[7:0]   ), //o
    .io_outputs_0_payload_counterDiff    (diffStage_controlPipe_fork_io_outputs_0_payload_counterDiff[7:0]), //o
    .io_outputs_0_payload_twiceCompValid (diffStage_controlPipe_fork_io_outputs_0_payload_twiceCompValid  ), //o
    .io_outputs_0_payload_twiceMode      (diffStage_controlPipe_fork_io_outputs_0_payload_twiceMode[2:0]  ), //o
    .io_outputs_1_valid                  (diffStage_controlPipe_fork_io_outputs_1_valid                   ), //o
    .io_outputs_1_ready                  (resultStage_pixelStream_ready                                   ), //i
    .io_outputs_1_payload_frameStart     (diffStage_controlPipe_fork_io_outputs_1_payload_frameStart      ), //o
    .io_outputs_1_payload_rowEnd         (diffStage_controlPipe_fork_io_outputs_1_payload_rowEnd          ), //o
    .io_outputs_1_payload_passMode       (diffStage_controlPipe_fork_io_outputs_1_payload_passMode        ), //o
    .io_outputs_1_payload_passValid      (diffStage_controlPipe_fork_io_outputs_1_payload_passValid       ), //o
    .io_outputs_1_payload_onceMode       (diffStage_controlPipe_fork_io_outputs_1_payload_onceMode[2:0]   ), //o
    .io_outputs_1_payload_onceValid      (diffStage_controlPipe_fork_io_outputs_1_payload_onceValid       ), //o
    .io_outputs_1_payload_mainCompare    (diffStage_controlPipe_fork_io_outputs_1_payload_mainCompare     ), //o
    .io_outputs_1_payload_counterCompare (diffStage_controlPipe_fork_io_outputs_1_payload_counterCompare  ), //o
    .io_outputs_1_payload_mainDiff       (diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff[7:0]   ), //o
    .io_outputs_1_payload_counterDiff    (diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff[7:0]), //o
    .io_outputs_1_payload_twiceCompValid (diffStage_controlPipe_fork_io_outputs_1_payload_twiceCompValid  ), //o
    .io_outputs_1_payload_twiceMode      (diffStage_controlPipe_fork_io_outputs_1_payload_twiceMode[2:0]  )  //o
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_BOOT : controlStateMachine_stateReg_string = "BOOT ";
      controlStateMachine_enumDef_HOLD : controlStateMachine_stateReg_string = "HOLD ";
      controlStateMachine_enumDef_PASS : controlStateMachine_stateReg_string = "PASS ";
      controlStateMachine_enumDef_ONCE : controlStateMachine_stateReg_string = "ONCE ";
      controlStateMachine_enumDef_TWICE : controlStateMachine_stateReg_string = "TWICE";
      default : controlStateMachine_stateReg_string = "?????";
    endcase
  end
  always @(*) begin
    case(controlStateMachine_stateNext)
      controlStateMachine_enumDef_BOOT : controlStateMachine_stateNext_string = "BOOT ";
      controlStateMachine_enumDef_HOLD : controlStateMachine_stateNext_string = "HOLD ";
      controlStateMachine_enumDef_PASS : controlStateMachine_stateNext_string = "PASS ";
      controlStateMachine_enumDef_ONCE : controlStateMachine_stateNext_string = "ONCE ";
      controlStateMachine_enumDef_TWICE : controlStateMachine_stateNext_string = "TWICE";
      default : controlStateMachine_stateNext_string = "?????";
    endcase
  end
  `endif

  always @(*) begin
    pixelsIn_ready = 1'b0;
    pixelsIn_ready = (! pixelsIn_rValid);
  end

  always @(*) begin
    pixelsOut_valid = 1'b0;
    pixelsOut_valid = pixelsStream_s2mPipe_m2sPipe_valid;
  end

  always @(*) begin
    pixelsOut_payload_pixel = 8'h0;
    pixelsOut_payload_pixel = pixelsStream_s2mPipe_m2sPipe_payload_pixel;
  end

  always @(*) begin
    pixelsOut_payload_frameStart = 1'b0;
    pixelsOut_payload_frameStart = pixelsStream_s2mPipe_m2sPipe_payload_frameStart;
  end

  always @(*) begin
    pixelsOut_payload_rowEnd = 1'b0;
    pixelsOut_payload_rowEnd = pixelsStream_s2mPipe_m2sPipe_payload_rowEnd;
  end

  always @(*) begin
    startOut = 1'b0;
    startOut = slaveStart;
  end

  always @(*) begin
    inpDoneOut = 1'b0;
    inpDoneOut = inpDone;
  end

  assign when_SuperResolutionPart1_l79 = (inpThreeDoneIn && inpTwoDoneIn);
  assign when_SuperResolutionPart1_l79_1 = (startIn && (! startIn_regNext));
  assign when_SuperResolutionPart1_l82 = (! startIn);
  assign when_SuperResolutionPart1_l85 = (startIn && (! readDone));
  assign when_SuperResolutionPart1_l85_1 = (! startIn);
  assign pixelsIn_fire = (pixelsIn_valid && pixelsIn_ready);
  assign when_SuperResolutionPart1_l88 = ((! inpTwoDoneIn) && pixelsIn_fire);
  assign when_SuperResolutionPart1_l88_1 = ((inpTwoDoneIn && inpThreeDoneIn) || (! startIn));
  assign when_SuperResolutionPart1_l103 = (! startIn);
  assign when_SuperResolutionPart1_l106 = (! startIn);
  always @(*) begin
    bufferRowCount_willIncrement = 1'b0;
    if(when_SuperResolutionPart1_l425) begin
      if(!bufferReachFinalRow) begin
        bufferRowCount_willIncrement = 1'b1;
      end
    end
  end

  always @(*) begin
    bufferRowCount_willClear = 1'b0;
    if(when_SuperResolutionPart1_l425) begin
      if(bufferReachFinalRow) begin
        bufferRowCount_willClear = 1'b1;
      end
    end
  end

  assign bufferRowCount_willOverflowIfInc = (bufferRowCount_value == 10'h21c);
  assign bufferRowCount_willOverflow = (bufferRowCount_willOverflowIfInc && bufferRowCount_willIncrement);
  always @(*) begin
    if(bufferRowCount_willOverflow) begin
      bufferRowCount_valueNext = 10'h0;
    end else begin
      bufferRowCount_valueNext = (bufferRowCount_value + CICC1851_bufferRowCount_valueNext);
    end
    if(bufferRowCount_willClear) begin
      bufferRowCount_valueNext = 10'h0;
    end
  end

  assign when_SuperResolutionPart1_l112 = ((startIn && (! holdBuffer)) && (! writeDone));
  assign when_SuperResolutionPart1_l112_1 = (((! startIn) || holdBuffer) || writeDone);
  assign when_SuperResolutionPart1_l115 = (! startRead);
  assign when_SuperResolutionPart1_l118 = (! startRead);
  always @(*) begin
    bufferWAddr_willIncrement = 1'b0;
    if(passPixels_fire_8) begin
      if(!passPixels_payload_rowEnd) begin
        bufferWAddr_willIncrement = 1'b1;
      end
    end
  end

  always @(*) begin
    bufferWAddr_willClear = 1'b0;
    if(passPixels_fire_8) begin
      if(passPixels_payload_rowEnd) begin
        bufferWAddr_willClear = 1'b1;
      end
    end
  end

  assign bufferWAddr_willOverflowIfInc = (bufferWAddr_value == 10'h3bf);
  assign bufferWAddr_willOverflow = (bufferWAddr_willOverflowIfInc && bufferWAddr_willIncrement);
  always @(*) begin
    if(bufferWAddr_willOverflow) begin
      bufferWAddr_valueNext = 10'h0;
    end else begin
      bufferWAddr_valueNext = (bufferWAddr_value + CICC1851_bufferWAddr_valueNext);
    end
    if(bufferWAddr_willClear) begin
      bufferWAddr_valueNext = 10'h0;
    end
  end

  always @(*) begin
    outPixelAddr_willIncrement = 1'b0;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_HOLD : begin
      end
      controlStateMachine_enumDef_PASS : begin
        if(controlStream_fire_6) begin
          if(!outReachRowEnd) begin
            outPixelAddr_willIncrement = 1'b1;
          end
        end
      end
      controlStateMachine_enumDef_ONCE : begin
        if(controlStream_fire_12) begin
          if(!outReachRowEnd) begin
            outPixelAddr_willIncrement = 1'b1;
          end
        end
      end
      controlStateMachine_enumDef_TWICE : begin
        if(controlStream_fire_17) begin
          if(!outReachRowEnd) begin
            outPixelAddr_willIncrement = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outPixelAddr_willClear = 1'b0;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_HOLD : begin
      end
      controlStateMachine_enumDef_PASS : begin
        if(controlStream_fire_6) begin
          if(outReachRowEnd) begin
            outPixelAddr_willClear = 1'b1;
          end
        end
      end
      controlStateMachine_enumDef_ONCE : begin
        if(controlStream_fire_12) begin
          if(outReachRowEnd) begin
            outPixelAddr_willClear = 1'b1;
          end
        end
      end
      controlStateMachine_enumDef_TWICE : begin
        if(controlStream_fire_17) begin
          if(outReachRowEnd) begin
            outPixelAddr_willClear = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign outPixelAddr_willOverflowIfInc = (outPixelAddr_value == 11'h77f);
  assign outPixelAddr_willOverflow = (outPixelAddr_willOverflowIfInc && outPixelAddr_willIncrement);
  always @(*) begin
    if(outPixelAddr_willOverflow) begin
      outPixelAddr_valueNext = 11'h0;
    end else begin
      outPixelAddr_valueNext = (outPixelAddr_value + CICC1851_outPixelAddr_valueNext);
    end
    if(outPixelAddr_willClear) begin
      outPixelAddr_valueNext = 11'h0;
    end
  end

  always @(*) begin
    outRowCount_willIncrement = 1'b0;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_HOLD : begin
      end
      controlStateMachine_enumDef_PASS : begin
        if(when_SuperResolutionPart1_l513) begin
          if(!outReachFinalRow) begin
            outRowCount_willIncrement = 1'b1;
          end
        end
      end
      controlStateMachine_enumDef_ONCE : begin
        if(when_SuperResolutionPart1_l581) begin
          if(!outReachFinalRow) begin
            outRowCount_willIncrement = 1'b1;
          end
        end
      end
      controlStateMachine_enumDef_TWICE : begin
        if(when_SuperResolutionPart1_l667) begin
          if(!outReachFinalRow) begin
            outRowCount_willIncrement = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outRowCount_willClear = 1'b0;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_HOLD : begin
      end
      controlStateMachine_enumDef_PASS : begin
        if(when_SuperResolutionPart1_l513) begin
          if(outReachFinalRow) begin
            outRowCount_willClear = 1'b1;
          end
        end
      end
      controlStateMachine_enumDef_ONCE : begin
        if(when_SuperResolutionPart1_l581) begin
          if(outReachFinalRow) begin
            outRowCount_willClear = 1'b1;
          end
        end
      end
      controlStateMachine_enumDef_TWICE : begin
        if(when_SuperResolutionPart1_l667) begin
          if(outReachFinalRow) begin
            outRowCount_willClear = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign outRowCount_willOverflowIfInc = (outRowCount_value == 11'h438);
  assign outRowCount_willOverflow = (outRowCount_willOverflowIfInc && outRowCount_willIncrement);
  always @(*) begin
    if(outRowCount_willOverflow) begin
      outRowCount_valueNext = 11'h0;
    end else begin
      outRowCount_valueNext = (outRowCount_value + CICC1851_outRowCount_valueNext);
    end
    if(outRowCount_willClear) begin
      outRowCount_valueNext = 11'h0;
    end
  end

  always @(*) begin
    mainAddrOne = CICC1851_mainAddrOne[9:0];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_HOLD : begin
      end
      controlStateMachine_enumDef_PASS : begin
      end
      controlStateMachine_enumDef_ONCE : begin
        if(when_SuperResolutionPart1_l537) begin
          if(nextRowBuffer) begin
            mainAddrOne = CICC1851_mainAddrOne_1[9:0];
          end
        end else begin
          mainAddrOne = CICC1851_mainAddrOne_3[9:0];
        end
      end
      controlStateMachine_enumDef_TWICE : begin
        if(outReachFinalRow) begin
          if(nextRowBuffer) begin
            if(outReachRowEnd) begin
              mainAddrOne = CICC1851_mainAddrOne_4[9:0];
            end else begin
              mainAddrOne = CICC1851_mainAddrOne_6[9:0];
            end
          end
        end else begin
          if(nextRowBuffer) begin
            mainAddrOne = CICC1851_mainAddrOne_8[9:0];
          end else begin
            if(outReachRowEnd) begin
              mainAddrOne = CICC1851_mainAddrOne_10[9:0];
            end else begin
              mainAddrOne = CICC1851_mainAddrOne_12[9:0];
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    counterAddrOne = CICC1851_counterAddrOne[9:0];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_HOLD : begin
      end
      controlStateMachine_enumDef_PASS : begin
      end
      controlStateMachine_enumDef_ONCE : begin
        if(when_SuperResolutionPart1_l537) begin
          if(nextRowBuffer) begin
            if(outReachRowEnd) begin
              counterAddrOne = CICC1851_counterAddrOne_1[9:0];
            end else begin
              counterAddrOne = CICC1851_counterAddrOne_3[9:0];
            end
          end
        end
      end
      controlStateMachine_enumDef_TWICE : begin
        if(outReachFinalRow) begin
          if(nextRowBuffer) begin
            if(!outReachRowEnd) begin
              counterAddrOne = CICC1851_counterAddrOne_7[9:0];
            end
          end
        end else begin
          if(nextRowBuffer) begin
            if(outReachRowEnd) begin
              counterAddrOne = CICC1851_counterAddrOne_11[9:0];
            end else begin
              counterAddrOne = CICC1851_counterAddrOne_13[9:0];
            end
          end else begin
            counterAddrOne = CICC1851_counterAddrOne_17[9:0];
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    mainAddrTwo = CICC1851_mainAddrTwo[9:0];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_HOLD : begin
      end
      controlStateMachine_enumDef_PASS : begin
      end
      controlStateMachine_enumDef_ONCE : begin
        if(when_SuperResolutionPart1_l537) begin
          if(!nextRowBuffer) begin
            mainAddrTwo = CICC1851_mainAddrTwo_1[9:0];
          end
        end else begin
          mainAddrTwo = CICC1851_mainAddrTwo_3[9:0];
        end
      end
      controlStateMachine_enumDef_TWICE : begin
        if(outReachFinalRow) begin
          if(!nextRowBuffer) begin
            if(outReachRowEnd) begin
              mainAddrTwo = CICC1851_mainAddrTwo_4[9:0];
            end else begin
              mainAddrTwo = CICC1851_mainAddrTwo_6[9:0];
            end
          end
        end else begin
          if(nextRowBuffer) begin
            if(outReachRowEnd) begin
              mainAddrTwo = CICC1851_mainAddrTwo_8[9:0];
            end else begin
              mainAddrTwo = CICC1851_mainAddrTwo_10[9:0];
            end
          end else begin
            mainAddrTwo = CICC1851_mainAddrTwo_14[9:0];
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    counterAddrTwo = CICC1851_counterAddrTwo[9:0];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_HOLD : begin
      end
      controlStateMachine_enumDef_PASS : begin
      end
      controlStateMachine_enumDef_ONCE : begin
        if(when_SuperResolutionPart1_l537) begin
          if(!nextRowBuffer) begin
            if(outReachRowEnd) begin
              counterAddrTwo = CICC1851_counterAddrTwo_1[9:0];
            end else begin
              counterAddrTwo = CICC1851_counterAddrTwo_3[9:0];
            end
          end
        end
      end
      controlStateMachine_enumDef_TWICE : begin
        if(outReachFinalRow) begin
          if(!nextRowBuffer) begin
            if(!outReachRowEnd) begin
              counterAddrTwo = CICC1851_counterAddrTwo_7[9:0];
            end
          end
        end else begin
          if(nextRowBuffer) begin
            counterAddrTwo = CICC1851_counterAddrTwo_11[9:0];
          end else begin
            if(outReachRowEnd) begin
              counterAddrTwo = CICC1851_counterAddrTwo_13[9:0];
            end else begin
              counterAddrTwo = CICC1851_counterAddrTwo_15[9:0];
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign validStream_valid = 1'b1;
  assign CICC1851_controls_frameStart = 30'h0;
  always @(*) begin
    controls_frameStart = CICC1851_controls_frameStart[0];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_HOLD : begin
      end
      controlStateMachine_enumDef_PASS : begin
        if(frameStart) begin
          controls_frameStart = 1'b1;
        end
      end
      controlStateMachine_enumDef_ONCE : begin
      end
      controlStateMachine_enumDef_TWICE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_rowEnd = CICC1851_controls_frameStart[1];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_HOLD : begin
      end
      controlStateMachine_enumDef_PASS : begin
        if(outReachRowEnd) begin
          controls_rowEnd = 1'b1;
        end
      end
      controlStateMachine_enumDef_ONCE : begin
        if(outReachRowEnd) begin
          controls_rowEnd = 1'b1;
        end
      end
      controlStateMachine_enumDef_TWICE : begin
        if(outReachRowEnd) begin
          controls_rowEnd = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_passMode = CICC1851_controls_frameStart[2];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_HOLD : begin
      end
      controlStateMachine_enumDef_PASS : begin
        if(nextRowBuffer) begin
          controls_passMode = 1'b0;
        end else begin
          controls_passMode = 1'b1;
        end
      end
      controlStateMachine_enumDef_ONCE : begin
      end
      controlStateMachine_enumDef_TWICE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_passValid = CICC1851_controls_frameStart[3];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_HOLD : begin
      end
      controlStateMachine_enumDef_PASS : begin
        controls_passValid = 1'b1;
      end
      controlStateMachine_enumDef_ONCE : begin
      end
      controlStateMachine_enumDef_TWICE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_onceMode = CICC1851_controls_frameStart[6 : 4];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_HOLD : begin
      end
      controlStateMachine_enumDef_PASS : begin
      end
      controlStateMachine_enumDef_ONCE : begin
        if(when_SuperResolutionPart1_l537) begin
          if(nextRowBuffer) begin
            controls_onceMode = 3'b000;
          end else begin
            controls_onceMode = {2'd0, CICC1851_controls_onceMode};
          end
        end else begin
          if(outReachFinalRow) begin
            if(nextRowBuffer) begin
              controls_onceMode = 3'b101;
            end else begin
              controls_onceMode = 3'b100;
            end
          end else begin
            if(nextRowBuffer) begin
              controls_onceMode = {1'd0, CICC1851_controls_onceMode_1};
            end else begin
              controls_onceMode = {1'd0, CICC1851_controls_onceMode_2};
            end
          end
        end
      end
      controlStateMachine_enumDef_TWICE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_onceValid = CICC1851_controls_frameStart[7];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_HOLD : begin
      end
      controlStateMachine_enumDef_PASS : begin
      end
      controlStateMachine_enumDef_ONCE : begin
        controls_onceValid = 1'b1;
      end
      controlStateMachine_enumDef_TWICE : begin
      end
      default : begin
      end
    endcase
  end

  assign controls_mainCompare = CICC1851_controls_frameStart[8];
  assign controls_counterCompare = CICC1851_controls_frameStart[9];
  assign controls_mainDiff = CICC1851_controls_frameStart[17 : 10];
  assign controls_counterDiff = CICC1851_controls_frameStart[25 : 18];
  always @(*) begin
    controls_twiceCompValid = CICC1851_controls_frameStart[26];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_HOLD : begin
      end
      controlStateMachine_enumDef_PASS : begin
      end
      controlStateMachine_enumDef_ONCE : begin
      end
      controlStateMachine_enumDef_TWICE : begin
        controls_twiceCompValid = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    controls_twiceMode = CICC1851_controls_frameStart[29 : 27];
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_HOLD : begin
      end
      controlStateMachine_enumDef_PASS : begin
      end
      controlStateMachine_enumDef_ONCE : begin
      end
      controlStateMachine_enumDef_TWICE : begin
        if(outReachFinalRow) begin
          if(nextRowBuffer) begin
            if(outReachRowEnd) begin
              controls_twiceMode = 3'b100;
            end else begin
              controls_twiceMode = 3'b101;
            end
          end else begin
            if(outReachRowEnd) begin
              controls_twiceMode = 3'b010;
            end else begin
              controls_twiceMode = 3'b011;
            end
          end
        end else begin
          if(nextRowBuffer) begin
            controls_twiceMode = 3'b000;
          end else begin
            controls_twiceMode = 3'b001;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    validStream_ready = (controlStream_ready && startRead);
    validStream_ready = (mainAddrOneStream_ready && startRead);
    validStream_ready = (counterAddrOneStream_ready && startRead);
    validStream_ready = (mainAddrTwoStream_ready && startRead);
    validStream_ready = (counterAddrTwoStream_ready && startRead);
  end

  assign controlStream_valid = (validStream_valid && startRead);
  assign controlStream_payload_frameStart = controls_frameStart;
  assign controlStream_payload_rowEnd = controls_rowEnd;
  assign controlStream_payload_passMode = controls_passMode;
  assign controlStream_payload_passValid = controls_passValid;
  assign controlStream_payload_onceMode = controls_onceMode;
  assign controlStream_payload_onceValid = controls_onceValid;
  assign controlStream_payload_mainCompare = controls_mainCompare;
  assign controlStream_payload_counterCompare = controls_counterCompare;
  assign controlStream_payload_mainDiff = controls_mainDiff;
  assign controlStream_payload_counterDiff = controls_counterDiff;
  assign controlStream_payload_twiceCompValid = controls_twiceCompValid;
  assign controlStream_payload_twiceMode = controls_twiceMode;
  assign mainAddrOneStream_valid = (validStream_valid && startRead);
  assign mainAddrOneStream_payload = mainAddrOne;
  assign counterAddrOneStream_valid = (validStream_valid && startRead);
  assign counterAddrOneStream_payload = counterAddrOne;
  assign mainAddrTwoStream_valid = (validStream_valid && startRead);
  assign mainAddrTwoStream_payload = mainAddrTwo;
  assign counterAddrTwoStream_valid = (validStream_valid && startRead);
  assign counterAddrTwoStream_payload = counterAddrTwo;
  assign mainAddrOneStream_ready = (! mainAddrOneStream_rValid);
  assign mainAddrOneStream_s2mPipe_valid = (mainAddrOneStream_valid || mainAddrOneStream_rValid);
  assign mainAddrOneStream_s2mPipe_payload = (mainAddrOneStream_rValid ? mainAddrOneStream_rData : mainAddrOneStream_payload);
  always @(*) begin
    mainAddrOneStream_s2mPipe_ready = mainAddrOneStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368) begin
      mainAddrOneStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368 = (! mainAddrOneStream_s2mPipe_m2sPipe_valid);
  assign mainAddrOneStream_s2mPipe_m2sPipe_valid = mainAddrOneStream_s2mPipe_rValid;
  assign mainAddrOneStream_s2mPipe_m2sPipe_payload = mainAddrOneStream_s2mPipe_rData;
  assign mainAddrOneStream_s2mPipe_m2sPipe_ready = ((! CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready) || CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready = CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_mainOnePixelStream_payload = CICC1851_lineBufferOne_port0;
  assign CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_1 = readStage_mainOnePixelStream_ready;
    if(when_Stream_l368_1) begin
      CICC1851_1 = 1'b1;
    end
  end

  assign when_Stream_l368_1 = (! readStage_mainOnePixelStream_valid);
  assign readStage_mainOnePixelStream_valid = CICC1851_readStage_mainOnePixelStream_valid;
  assign readStage_mainOnePixelStream_payload = CICC1851_readStage_mainOnePixelStream_payload_2;
  assign counterAddrOneStream_ready = (! counterAddrOneStream_rValid);
  assign counterAddrOneStream_s2mPipe_valid = (counterAddrOneStream_valid || counterAddrOneStream_rValid);
  assign counterAddrOneStream_s2mPipe_payload = (counterAddrOneStream_rValid ? counterAddrOneStream_rData : counterAddrOneStream_payload);
  always @(*) begin
    counterAddrOneStream_s2mPipe_ready = counterAddrOneStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_2) begin
      counterAddrOneStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_2 = (! counterAddrOneStream_s2mPipe_m2sPipe_valid);
  assign counterAddrOneStream_s2mPipe_m2sPipe_valid = counterAddrOneStream_s2mPipe_rValid;
  assign counterAddrOneStream_s2mPipe_m2sPipe_payload = counterAddrOneStream_s2mPipe_rData;
  assign counterAddrOneStream_s2mPipe_m2sPipe_ready = ((! CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready) || CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready = CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_counterOnePixelStream_payload = CICC1851_lineBufferOne_port1;
  assign CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_2 = readStage_counterOnePixelStream_ready;
    if(when_Stream_l368_3) begin
      CICC1851_2 = 1'b1;
    end
  end

  assign when_Stream_l368_3 = (! readStage_counterOnePixelStream_valid);
  assign readStage_counterOnePixelStream_valid = CICC1851_readStage_counterOnePixelStream_valid;
  assign readStage_counterOnePixelStream_payload = CICC1851_readStage_counterOnePixelStream_payload_2;
  assign mainAddrTwoStream_ready = (! mainAddrTwoStream_rValid);
  assign mainAddrTwoStream_s2mPipe_valid = (mainAddrTwoStream_valid || mainAddrTwoStream_rValid);
  assign mainAddrTwoStream_s2mPipe_payload = (mainAddrTwoStream_rValid ? mainAddrTwoStream_rData : mainAddrTwoStream_payload);
  always @(*) begin
    mainAddrTwoStream_s2mPipe_ready = mainAddrTwoStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_4) begin
      mainAddrTwoStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_4 = (! mainAddrTwoStream_s2mPipe_m2sPipe_valid);
  assign mainAddrTwoStream_s2mPipe_m2sPipe_valid = mainAddrTwoStream_s2mPipe_rValid;
  assign mainAddrTwoStream_s2mPipe_m2sPipe_payload = mainAddrTwoStream_s2mPipe_rData;
  assign mainAddrTwoStream_s2mPipe_m2sPipe_ready = ((! CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready) || CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready = CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_mainTwoPixelStream_payload = CICC1851_lineBufferTwo_port0;
  assign CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_3 = readStage_mainTwoPixelStream_ready;
    if(when_Stream_l368_5) begin
      CICC1851_3 = 1'b1;
    end
  end

  assign when_Stream_l368_5 = (! readStage_mainTwoPixelStream_valid);
  assign readStage_mainTwoPixelStream_valid = CICC1851_readStage_mainTwoPixelStream_valid;
  assign readStage_mainTwoPixelStream_payload = CICC1851_readStage_mainTwoPixelStream_payload_2;
  assign counterAddrTwoStream_ready = (! counterAddrTwoStream_rValid);
  assign counterAddrTwoStream_s2mPipe_valid = (counterAddrTwoStream_valid || counterAddrTwoStream_rValid);
  assign counterAddrTwoStream_s2mPipe_payload = (counterAddrTwoStream_rValid ? counterAddrTwoStream_rData : counterAddrTwoStream_payload);
  always @(*) begin
    counterAddrTwoStream_s2mPipe_ready = counterAddrTwoStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_6) begin
      counterAddrTwoStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_6 = (! counterAddrTwoStream_s2mPipe_m2sPipe_valid);
  assign counterAddrTwoStream_s2mPipe_m2sPipe_valid = counterAddrTwoStream_s2mPipe_rValid;
  assign counterAddrTwoStream_s2mPipe_m2sPipe_payload = counterAddrTwoStream_s2mPipe_rData;
  assign counterAddrTwoStream_s2mPipe_m2sPipe_ready = ((! CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready) || CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_1);
  assign CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready = CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_2;
  assign CICC1851_readStage_counterTwoPixelStream_payload = CICC1851_lineBufferTwo_port1;
  assign CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_1 = (! CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_3);
  always @(*) begin
    CICC1851_4 = readStage_counterTwoPixelStream_ready;
    if(when_Stream_l368_7) begin
      CICC1851_4 = 1'b1;
    end
  end

  assign when_Stream_l368_7 = (! readStage_counterTwoPixelStream_valid);
  assign readStage_counterTwoPixelStream_valid = CICC1851_readStage_counterTwoPixelStream_valid;
  assign readStage_counterTwoPixelStream_payload = CICC1851_readStage_counterTwoPixelStream_payload_2;
  assign controlStream_ready = (! controlStream_rValid);
  assign controlStream_s2mPipe_valid = (controlStream_valid || controlStream_rValid);
  assign controlStream_s2mPipe_payload_frameStart = (controlStream_rValid ? controlStream_rData_frameStart : controlStream_payload_frameStart);
  assign controlStream_s2mPipe_payload_rowEnd = (controlStream_rValid ? controlStream_rData_rowEnd : controlStream_payload_rowEnd);
  assign controlStream_s2mPipe_payload_passMode = (controlStream_rValid ? controlStream_rData_passMode : controlStream_payload_passMode);
  assign controlStream_s2mPipe_payload_passValid = (controlStream_rValid ? controlStream_rData_passValid : controlStream_payload_passValid);
  assign controlStream_s2mPipe_payload_onceMode = (controlStream_rValid ? controlStream_rData_onceMode : controlStream_payload_onceMode);
  assign controlStream_s2mPipe_payload_onceValid = (controlStream_rValid ? controlStream_rData_onceValid : controlStream_payload_onceValid);
  assign controlStream_s2mPipe_payload_mainCompare = (controlStream_rValid ? controlStream_rData_mainCompare : controlStream_payload_mainCompare);
  assign controlStream_s2mPipe_payload_counterCompare = (controlStream_rValid ? controlStream_rData_counterCompare : controlStream_payload_counterCompare);
  assign controlStream_s2mPipe_payload_mainDiff = (controlStream_rValid ? controlStream_rData_mainDiff : controlStream_payload_mainDiff);
  assign controlStream_s2mPipe_payload_counterDiff = (controlStream_rValid ? controlStream_rData_counterDiff : controlStream_payload_counterDiff);
  assign controlStream_s2mPipe_payload_twiceCompValid = (controlStream_rValid ? controlStream_rData_twiceCompValid : controlStream_payload_twiceCompValid);
  assign controlStream_s2mPipe_payload_twiceMode = (controlStream_rValid ? controlStream_rData_twiceMode : controlStream_payload_twiceMode);
  always @(*) begin
    controlStream_s2mPipe_ready = controlStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_8) begin
      controlStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_8 = (! controlStream_s2mPipe_m2sPipe_valid);
  assign controlStream_s2mPipe_m2sPipe_valid = controlStream_s2mPipe_rValid;
  assign controlStream_s2mPipe_m2sPipe_payload_frameStart = controlStream_s2mPipe_rData_frameStart;
  assign controlStream_s2mPipe_m2sPipe_payload_rowEnd = controlStream_s2mPipe_rData_rowEnd;
  assign controlStream_s2mPipe_m2sPipe_payload_passMode = controlStream_s2mPipe_rData_passMode;
  assign controlStream_s2mPipe_m2sPipe_payload_passValid = controlStream_s2mPipe_rData_passValid;
  assign controlStream_s2mPipe_m2sPipe_payload_onceMode = controlStream_s2mPipe_rData_onceMode;
  assign controlStream_s2mPipe_m2sPipe_payload_onceValid = controlStream_s2mPipe_rData_onceValid;
  assign controlStream_s2mPipe_m2sPipe_payload_mainCompare = controlStream_s2mPipe_rData_mainCompare;
  assign controlStream_s2mPipe_m2sPipe_payload_counterCompare = controlStream_s2mPipe_rData_counterCompare;
  assign controlStream_s2mPipe_m2sPipe_payload_mainDiff = controlStream_s2mPipe_rData_mainDiff;
  assign controlStream_s2mPipe_m2sPipe_payload_counterDiff = controlStream_s2mPipe_rData_counterDiff;
  assign controlStream_s2mPipe_m2sPipe_payload_twiceCompValid = controlStream_s2mPipe_rData_twiceCompValid;
  assign controlStream_s2mPipe_m2sPipe_payload_twiceMode = controlStream_s2mPipe_rData_twiceMode;
  always @(*) begin
    controlStream_s2mPipe_m2sPipe_ready = controlStream_s2mPipe_m2sPipe_m2sPipe_ready;
    if(when_Stream_l368_9) begin
      controlStream_s2mPipe_m2sPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_9 = (! controlStream_s2mPipe_m2sPipe_m2sPipe_valid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_valid = controlStream_s2mPipe_m2sPipe_rValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_frameStart = controlStream_s2mPipe_m2sPipe_rData_frameStart;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_rowEnd = controlStream_s2mPipe_m2sPipe_rData_rowEnd;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passMode = controlStream_s2mPipe_m2sPipe_rData_passMode;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passValid = controlStream_s2mPipe_m2sPipe_rData_passValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceMode = controlStream_s2mPipe_m2sPipe_rData_onceMode;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceValid = controlStream_s2mPipe_m2sPipe_rData_onceValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainCompare = controlStream_s2mPipe_m2sPipe_rData_mainCompare;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterCompare = controlStream_s2mPipe_m2sPipe_rData_counterCompare;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDiff = controlStream_s2mPipe_m2sPipe_rData_mainDiff;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDiff = controlStream_s2mPipe_m2sPipe_rData_counterDiff;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceCompValid = controlStream_s2mPipe_m2sPipe_rData_twiceCompValid;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceMode = controlStream_s2mPipe_m2sPipe_rData_twiceMode;
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_ready = (! controlStream_s2mPipe_m2sPipe_m2sPipe_rValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_valid = (controlStream_s2mPipe_m2sPipe_m2sPipe_valid || controlStream_s2mPipe_m2sPipe_m2sPipe_rValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_frameStart = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_frameStart : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_frameStart);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_rowEnd = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_rowEnd : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_rowEnd);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_passMode = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_passMode : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passMode);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_passValid = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_passValid : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_onceMode = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_onceMode : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceMode);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_onceValid = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_onceValid : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainCompare = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainCompare : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainCompare);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterCompare = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterCompare : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterCompare);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainDiff = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainDiff : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDiff);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterDiff = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterDiff : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDiff);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_twiceCompValid = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_twiceCompValid : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceCompValid);
  assign controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_twiceMode = (controlStream_s2mPipe_m2sPipe_m2sPipe_rValid ? controlStream_s2mPipe_m2sPipe_m2sPipe_rData_twiceMode : controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceMode);
  always @(*) begin
    controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready = readStage_controlPipe_ready;
    if(when_Stream_l368_10) begin
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_10 = (! readStage_controlPipe_valid);
  assign readStage_controlPipe_valid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rValid;
  assign readStage_controlPipe_payload_frameStart = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_frameStart;
  assign readStage_controlPipe_payload_rowEnd = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_rowEnd;
  assign readStage_controlPipe_payload_passMode = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_passMode;
  assign readStage_controlPipe_payload_passValid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_passValid;
  assign readStage_controlPipe_payload_onceMode = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_onceMode;
  assign readStage_controlPipe_payload_onceValid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_onceValid;
  assign readStage_controlPipe_payload_mainCompare = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainCompare;
  assign readStage_controlPipe_payload_counterCompare = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterCompare;
  assign readStage_controlPipe_payload_mainDiff = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainDiff;
  assign readStage_controlPipe_payload_counterDiff = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterDiff;
  assign readStage_controlPipe_payload_twiceCompValid = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_twiceCompValid;
  assign readStage_controlPipe_payload_twiceMode = controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_twiceMode;
  assign readStage_mainOnePixelStream_ready = (! readStage_mainOnePixelStream_rValid);
  assign readStage_mainOnePixelStream_s2mPipe_valid = (readStage_mainOnePixelStream_valid || readStage_mainOnePixelStream_rValid);
  assign readStage_mainOnePixelStream_s2mPipe_payload = (readStage_mainOnePixelStream_rValid ? readStage_mainOnePixelStream_rData : readStage_mainOnePixelStream_payload);
  always @(*) begin
    readStage_mainOnePixelStream_s2mPipe_ready = compareStage_mainOnePixelStream_ready;
    if(when_Stream_l368_11) begin
      readStage_mainOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_11 = (! compareStage_mainOnePixelStream_valid);
  assign compareStage_mainOnePixelStream_valid = readStage_mainOnePixelStream_s2mPipe_rValid;
  assign compareStage_mainOnePixelStream_payload = readStage_mainOnePixelStream_s2mPipe_rData;
  assign readStage_counterOnePixelStream_ready = (! readStage_counterOnePixelStream_rValid);
  assign readStage_counterOnePixelStream_s2mPipe_valid = (readStage_counterOnePixelStream_valid || readStage_counterOnePixelStream_rValid);
  assign readStage_counterOnePixelStream_s2mPipe_payload = (readStage_counterOnePixelStream_rValid ? readStage_counterOnePixelStream_rData : readStage_counterOnePixelStream_payload);
  always @(*) begin
    readStage_counterOnePixelStream_s2mPipe_ready = compareStage_counterOnePixelStream_ready;
    if(when_Stream_l368_12) begin
      readStage_counterOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_12 = (! compareStage_counterOnePixelStream_valid);
  assign compareStage_counterOnePixelStream_valid = readStage_counterOnePixelStream_s2mPipe_rValid;
  assign compareStage_counterOnePixelStream_payload = readStage_counterOnePixelStream_s2mPipe_rData;
  assign readStage_mainTwoPixelStream_ready = (! readStage_mainTwoPixelStream_rValid);
  assign readStage_mainTwoPixelStream_s2mPipe_valid = (readStage_mainTwoPixelStream_valid || readStage_mainTwoPixelStream_rValid);
  assign readStage_mainTwoPixelStream_s2mPipe_payload = (readStage_mainTwoPixelStream_rValid ? readStage_mainTwoPixelStream_rData : readStage_mainTwoPixelStream_payload);
  always @(*) begin
    readStage_mainTwoPixelStream_s2mPipe_ready = compareStage_mainTwoPixelStream_ready;
    if(when_Stream_l368_13) begin
      readStage_mainTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_13 = (! compareStage_mainTwoPixelStream_valid);
  assign compareStage_mainTwoPixelStream_valid = readStage_mainTwoPixelStream_s2mPipe_rValid;
  assign compareStage_mainTwoPixelStream_payload = readStage_mainTwoPixelStream_s2mPipe_rData;
  assign readStage_counterTwoPixelStream_ready = (! readStage_counterTwoPixelStream_rValid);
  assign readStage_counterTwoPixelStream_s2mPipe_valid = (readStage_counterTwoPixelStream_valid || readStage_counterTwoPixelStream_rValid);
  assign readStage_counterTwoPixelStream_s2mPipe_payload = (readStage_counterTwoPixelStream_rValid ? readStage_counterTwoPixelStream_rData : readStage_counterTwoPixelStream_payload);
  always @(*) begin
    readStage_counterTwoPixelStream_s2mPipe_ready = compareStage_counterTwoPixelStream_ready;
    if(when_Stream_l368_14) begin
      readStage_counterTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_14 = (! compareStage_counterTwoPixelStream_valid);
  assign compareStage_counterTwoPixelStream_valid = readStage_counterTwoPixelStream_s2mPipe_rValid;
  assign compareStage_counterTwoPixelStream_payload = readStage_counterTwoPixelStream_s2mPipe_rData;
  always @(*) begin
    CICC1851_readStage_controlPipe_translated_payload_mainCompare = readStage_controlPipe_payload_mainCompare;
    if(readStage_controlPipe_payload_onceValid) begin
      case(readStage_controlPipe_payload_onceMode)
        3'b000 : begin
          if(when_SuperResolutionPart1_l205) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        3'b001 : begin
          if(when_SuperResolutionPart1_l209) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        3'b010 : begin
          if(when_SuperResolutionPart1_l213) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        3'b011 : begin
          if(when_SuperResolutionPart1_l217) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        3'b100 : begin
          CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
        end
        3'b101 : begin
          CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
        end
        default : begin
        end
      endcase
    end
    if(readStage_controlPipe_payload_twiceCompValid) begin
      case(readStage_controlPipe_payload_twiceMode)
        3'b000 : begin
          if(when_SuperResolutionPart1_l228) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        3'b001 : begin
          if(when_SuperResolutionPart1_l234) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        3'b010 : begin
          CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
        end
        3'b011 : begin
          if(when_SuperResolutionPart1_l241) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        3'b100 : begin
          CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
        end
        3'b101 : begin
          if(when_SuperResolutionPart1_l246) begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_mainCompare = 1'b0;
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    CICC1851_readStage_controlPipe_translated_payload_counterCompare = readStage_controlPipe_payload_counterCompare;
    if(readStage_controlPipe_payload_twiceCompValid) begin
      case(readStage_controlPipe_payload_twiceMode)
        3'b000 : begin
          if(when_SuperResolutionPart1_l230) begin
            CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
          end
        end
        3'b001 : begin
          if(when_SuperResolutionPart1_l236) begin
            CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b1;
          end else begin
            CICC1851_readStage_controlPipe_translated_payload_counterCompare = 1'b0;
          end
        end
        default : begin
        end
      endcase
    end
  end

  assign when_SuperResolutionPart1_l205 = (readStage_counterOnePixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart1_l209 = (readStage_counterTwoPixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart1_l213 = (readStage_mainTwoPixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart1_l217 = (readStage_mainOnePixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart1_l228 = (readStage_mainTwoPixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign when_SuperResolutionPart1_l230 = (readStage_counterOnePixelStream_payload <= readStage_counterTwoPixelStream_payload);
  assign when_SuperResolutionPart1_l234 = (readStage_mainOnePixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart1_l236 = (readStage_counterTwoPixelStream_payload <= readStage_counterOnePixelStream_payload);
  assign when_SuperResolutionPart1_l241 = (readStage_counterTwoPixelStream_payload <= readStage_mainTwoPixelStream_payload);
  assign when_SuperResolutionPart1_l246 = (readStage_counterOnePixelStream_payload <= readStage_mainOnePixelStream_payload);
  assign readStage_controlPipe_translated_valid = readStage_controlPipe_valid;
  assign readStage_controlPipe_ready = readStage_controlPipe_translated_ready;
  assign readStage_controlPipe_translated_payload_frameStart = readStage_controlPipe_payload_frameStart;
  assign readStage_controlPipe_translated_payload_rowEnd = readStage_controlPipe_payload_rowEnd;
  assign readStage_controlPipe_translated_payload_passMode = readStage_controlPipe_payload_passMode;
  assign readStage_controlPipe_translated_payload_passValid = readStage_controlPipe_payload_passValid;
  assign readStage_controlPipe_translated_payload_onceMode = readStage_controlPipe_payload_onceMode;
  assign readStage_controlPipe_translated_payload_onceValid = readStage_controlPipe_payload_onceValid;
  assign readStage_controlPipe_translated_payload_mainCompare = CICC1851_readStage_controlPipe_translated_payload_mainCompare;
  assign readStage_controlPipe_translated_payload_counterCompare = CICC1851_readStage_controlPipe_translated_payload_counterCompare;
  assign readStage_controlPipe_translated_payload_mainDiff = readStage_controlPipe_payload_mainDiff;
  assign readStage_controlPipe_translated_payload_counterDiff = readStage_controlPipe_payload_counterDiff;
  assign readStage_controlPipe_translated_payload_twiceCompValid = readStage_controlPipe_payload_twiceCompValid;
  assign readStage_controlPipe_translated_payload_twiceMode = readStage_controlPipe_payload_twiceMode;
  assign readStage_controlPipe_translated_ready = (! readStage_controlPipe_translated_rValid);
  assign readStage_controlPipe_translated_s2mPipe_valid = (readStage_controlPipe_translated_valid || readStage_controlPipe_translated_rValid);
  assign readStage_controlPipe_translated_s2mPipe_payload_frameStart = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_frameStart : readStage_controlPipe_translated_payload_frameStart);
  assign readStage_controlPipe_translated_s2mPipe_payload_rowEnd = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_rowEnd : readStage_controlPipe_translated_payload_rowEnd);
  assign readStage_controlPipe_translated_s2mPipe_payload_passMode = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_passMode : readStage_controlPipe_translated_payload_passMode);
  assign readStage_controlPipe_translated_s2mPipe_payload_passValid = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_passValid : readStage_controlPipe_translated_payload_passValid);
  assign readStage_controlPipe_translated_s2mPipe_payload_onceMode = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_onceMode : readStage_controlPipe_translated_payload_onceMode);
  assign readStage_controlPipe_translated_s2mPipe_payload_onceValid = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_onceValid : readStage_controlPipe_translated_payload_onceValid);
  assign readStage_controlPipe_translated_s2mPipe_payload_mainCompare = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_mainCompare : readStage_controlPipe_translated_payload_mainCompare);
  assign readStage_controlPipe_translated_s2mPipe_payload_counterCompare = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_counterCompare : readStage_controlPipe_translated_payload_counterCompare);
  assign readStage_controlPipe_translated_s2mPipe_payload_mainDiff = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_mainDiff : readStage_controlPipe_translated_payload_mainDiff);
  assign readStage_controlPipe_translated_s2mPipe_payload_counterDiff = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_counterDiff : readStage_controlPipe_translated_payload_counterDiff);
  assign readStage_controlPipe_translated_s2mPipe_payload_twiceCompValid = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_twiceCompValid : readStage_controlPipe_translated_payload_twiceCompValid);
  assign readStage_controlPipe_translated_s2mPipe_payload_twiceMode = (readStage_controlPipe_translated_rValid ? readStage_controlPipe_translated_rData_twiceMode : readStage_controlPipe_translated_payload_twiceMode);
  always @(*) begin
    readStage_controlPipe_translated_s2mPipe_ready = compareStage_controlPipe_ready;
    if(when_Stream_l368_15) begin
      readStage_controlPipe_translated_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_15 = (! compareStage_controlPipe_valid);
  assign compareStage_controlPipe_valid = readStage_controlPipe_translated_s2mPipe_rValid;
  assign compareStage_controlPipe_payload_frameStart = readStage_controlPipe_translated_s2mPipe_rData_frameStart;
  assign compareStage_controlPipe_payload_rowEnd = readStage_controlPipe_translated_s2mPipe_rData_rowEnd;
  assign compareStage_controlPipe_payload_passMode = readStage_controlPipe_translated_s2mPipe_rData_passMode;
  assign compareStage_controlPipe_payload_passValid = readStage_controlPipe_translated_s2mPipe_rData_passValid;
  assign compareStage_controlPipe_payload_onceMode = readStage_controlPipe_translated_s2mPipe_rData_onceMode;
  assign compareStage_controlPipe_payload_onceValid = readStage_controlPipe_translated_s2mPipe_rData_onceValid;
  assign compareStage_controlPipe_payload_mainCompare = readStage_controlPipe_translated_s2mPipe_rData_mainCompare;
  assign compareStage_controlPipe_payload_counterCompare = readStage_controlPipe_translated_s2mPipe_rData_counterCompare;
  assign compareStage_controlPipe_payload_mainDiff = readStage_controlPipe_translated_s2mPipe_rData_mainDiff;
  assign compareStage_controlPipe_payload_counterDiff = readStage_controlPipe_translated_s2mPipe_rData_counterDiff;
  assign compareStage_controlPipe_payload_twiceCompValid = readStage_controlPipe_translated_s2mPipe_rData_twiceCompValid;
  assign compareStage_controlPipe_payload_twiceMode = readStage_controlPipe_translated_s2mPipe_rData_twiceMode;
  assign compareStage_mainOnePixelStream_ready = (! compareStage_mainOnePixelStream_rValid);
  assign compareStage_mainOnePixelStream_s2mPipe_valid = (compareStage_mainOnePixelStream_valid || compareStage_mainOnePixelStream_rValid);
  assign compareStage_mainOnePixelStream_s2mPipe_payload = (compareStage_mainOnePixelStream_rValid ? compareStage_mainOnePixelStream_rData : compareStage_mainOnePixelStream_payload);
  always @(*) begin
    compareStage_mainOnePixelStream_s2mPipe_ready = diffStage_mainOnePixelStream_ready;
    if(when_Stream_l368_16) begin
      compareStage_mainOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_16 = (! diffStage_mainOnePixelStream_valid);
  assign diffStage_mainOnePixelStream_valid = compareStage_mainOnePixelStream_s2mPipe_rValid;
  assign diffStage_mainOnePixelStream_payload = compareStage_mainOnePixelStream_s2mPipe_rData;
  assign compareStage_counterOnePixelStream_ready = (! compareStage_counterOnePixelStream_rValid);
  assign compareStage_counterOnePixelStream_s2mPipe_valid = (compareStage_counterOnePixelStream_valid || compareStage_counterOnePixelStream_rValid);
  assign compareStage_counterOnePixelStream_s2mPipe_payload = (compareStage_counterOnePixelStream_rValid ? compareStage_counterOnePixelStream_rData : compareStage_counterOnePixelStream_payload);
  always @(*) begin
    compareStage_counterOnePixelStream_s2mPipe_ready = diffStage_counterOnePixelStream_ready;
    if(when_Stream_l368_17) begin
      compareStage_counterOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_17 = (! diffStage_counterOnePixelStream_valid);
  assign diffStage_counterOnePixelStream_valid = compareStage_counterOnePixelStream_s2mPipe_rValid;
  assign diffStage_counterOnePixelStream_payload = compareStage_counterOnePixelStream_s2mPipe_rData;
  assign compareStage_mainTwoPixelStream_ready = (! compareStage_mainTwoPixelStream_rValid);
  assign compareStage_mainTwoPixelStream_s2mPipe_valid = (compareStage_mainTwoPixelStream_valid || compareStage_mainTwoPixelStream_rValid);
  assign compareStage_mainTwoPixelStream_s2mPipe_payload = (compareStage_mainTwoPixelStream_rValid ? compareStage_mainTwoPixelStream_rData : compareStage_mainTwoPixelStream_payload);
  always @(*) begin
    compareStage_mainTwoPixelStream_s2mPipe_ready = diffStage_mainTwoPixelStream_ready;
    if(when_Stream_l368_18) begin
      compareStage_mainTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_18 = (! diffStage_mainTwoPixelStream_valid);
  assign diffStage_mainTwoPixelStream_valid = compareStage_mainTwoPixelStream_s2mPipe_rValid;
  assign diffStage_mainTwoPixelStream_payload = compareStage_mainTwoPixelStream_s2mPipe_rData;
  assign compareStage_counterTwoPixelStream_ready = (! compareStage_counterTwoPixelStream_rValid);
  assign compareStage_counterTwoPixelStream_s2mPipe_valid = (compareStage_counterTwoPixelStream_valid || compareStage_counterTwoPixelStream_rValid);
  assign compareStage_counterTwoPixelStream_s2mPipe_payload = (compareStage_counterTwoPixelStream_rValid ? compareStage_counterTwoPixelStream_rData : compareStage_counterTwoPixelStream_payload);
  always @(*) begin
    compareStage_counterTwoPixelStream_s2mPipe_ready = diffStage_counterTwoPixelStream_ready;
    if(when_Stream_l368_19) begin
      compareStage_counterTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_19 = (! diffStage_counterTwoPixelStream_valid);
  assign diffStage_counterTwoPixelStream_valid = compareStage_counterTwoPixelStream_s2mPipe_rValid;
  assign diffStage_counterTwoPixelStream_payload = compareStage_counterTwoPixelStream_s2mPipe_rData;
  always @(*) begin
    CICC1851_compareStage_controlPipe_translated_payload_mainDiff = compareStage_controlPipe_payload_mainDiff;
    if(compareStage_controlPipe_payload_onceValid) begin
      case(compareStage_controlPipe_payload_onceMode)
        3'b000 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_counterOnePixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterOnePixelStream_payload - compareStage_mainOnePixelStream_payload);
          end
        end
        3'b001 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterTwoPixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainTwoPixelStream_payload);
          end
        end
        3'b010 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_mainTwoPixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_mainOnePixelStream_payload);
          end
        end
        3'b011 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_mainOnePixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_mainTwoPixelStream_payload);
          end
        end
        3'b100 : begin
          CICC1851_compareStage_controlPipe_translated_payload_mainDiff = 8'h0;
        end
        3'b101 : begin
          CICC1851_compareStage_controlPipe_translated_payload_mainDiff = 8'h0;
        end
        default : begin
        end
      endcase
    end
    if(compareStage_controlPipe_payload_twiceCompValid) begin
      case(compareStage_controlPipe_payload_twiceMode)
        3'b000 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_mainTwoPixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_mainOnePixelStream_payload);
          end
        end
        3'b001 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_mainOnePixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_mainTwoPixelStream_payload);
          end
        end
        3'b010 : begin
          CICC1851_compareStage_controlPipe_translated_payload_mainDiff = 8'h0;
        end
        3'b011 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainTwoPixelStream_payload - compareStage_counterTwoPixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterTwoPixelStream_payload - compareStage_mainTwoPixelStream_payload);
          end
        end
        3'b100 : begin
          CICC1851_compareStage_controlPipe_translated_payload_mainDiff = 8'h0;
        end
        3'b101 : begin
          if(compareStage_controlPipe_payload_mainCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_mainOnePixelStream_payload - compareStage_counterOnePixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_mainDiff = (compareStage_counterOnePixelStream_payload - compareStage_mainOnePixelStream_payload);
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    CICC1851_compareStage_controlPipe_translated_payload_counterDiff = compareStage_controlPipe_payload_counterDiff;
    if(compareStage_controlPipe_payload_twiceCompValid) begin
      case(compareStage_controlPipe_payload_twiceMode)
        3'b000 : begin
          if(compareStage_controlPipe_payload_counterCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterTwoPixelStream_payload - compareStage_counterOnePixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterOnePixelStream_payload - compareStage_counterTwoPixelStream_payload);
          end
        end
        3'b001 : begin
          if(compareStage_controlPipe_payload_counterCompare) begin
            CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterOnePixelStream_payload - compareStage_counterTwoPixelStream_payload);
          end else begin
            CICC1851_compareStage_controlPipe_translated_payload_counterDiff = (compareStage_counterTwoPixelStream_payload - compareStage_counterOnePixelStream_payload);
          end
        end
        default : begin
        end
      endcase
    end
  end

  assign compareStage_controlPipe_translated_valid = compareStage_controlPipe_valid;
  assign compareStage_controlPipe_ready = compareStage_controlPipe_translated_ready;
  assign compareStage_controlPipe_translated_payload_frameStart = compareStage_controlPipe_payload_frameStart;
  assign compareStage_controlPipe_translated_payload_rowEnd = compareStage_controlPipe_payload_rowEnd;
  assign compareStage_controlPipe_translated_payload_passMode = compareStage_controlPipe_payload_passMode;
  assign compareStage_controlPipe_translated_payload_passValid = compareStage_controlPipe_payload_passValid;
  assign compareStage_controlPipe_translated_payload_onceMode = compareStage_controlPipe_payload_onceMode;
  assign compareStage_controlPipe_translated_payload_onceValid = compareStage_controlPipe_payload_onceValid;
  assign compareStage_controlPipe_translated_payload_mainCompare = compareStage_controlPipe_payload_mainCompare;
  assign compareStage_controlPipe_translated_payload_counterCompare = compareStage_controlPipe_payload_counterCompare;
  assign compareStage_controlPipe_translated_payload_mainDiff = CICC1851_compareStage_controlPipe_translated_payload_mainDiff;
  assign compareStage_controlPipe_translated_payload_counterDiff = CICC1851_compareStage_controlPipe_translated_payload_counterDiff;
  assign compareStage_controlPipe_translated_payload_twiceCompValid = compareStage_controlPipe_payload_twiceCompValid;
  assign compareStage_controlPipe_translated_payload_twiceMode = compareStage_controlPipe_payload_twiceMode;
  assign compareStage_controlPipe_translated_ready = (! compareStage_controlPipe_translated_rValid);
  assign compareStage_controlPipe_translated_s2mPipe_valid = (compareStage_controlPipe_translated_valid || compareStage_controlPipe_translated_rValid);
  assign compareStage_controlPipe_translated_s2mPipe_payload_frameStart = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_frameStart : compareStage_controlPipe_translated_payload_frameStart);
  assign compareStage_controlPipe_translated_s2mPipe_payload_rowEnd = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_rowEnd : compareStage_controlPipe_translated_payload_rowEnd);
  assign compareStage_controlPipe_translated_s2mPipe_payload_passMode = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_passMode : compareStage_controlPipe_translated_payload_passMode);
  assign compareStage_controlPipe_translated_s2mPipe_payload_passValid = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_passValid : compareStage_controlPipe_translated_payload_passValid);
  assign compareStage_controlPipe_translated_s2mPipe_payload_onceMode = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_onceMode : compareStage_controlPipe_translated_payload_onceMode);
  assign compareStage_controlPipe_translated_s2mPipe_payload_onceValid = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_onceValid : compareStage_controlPipe_translated_payload_onceValid);
  assign compareStage_controlPipe_translated_s2mPipe_payload_mainCompare = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_mainCompare : compareStage_controlPipe_translated_payload_mainCompare);
  assign compareStage_controlPipe_translated_s2mPipe_payload_counterCompare = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_counterCompare : compareStage_controlPipe_translated_payload_counterCompare);
  assign compareStage_controlPipe_translated_s2mPipe_payload_mainDiff = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_mainDiff : compareStage_controlPipe_translated_payload_mainDiff);
  assign compareStage_controlPipe_translated_s2mPipe_payload_counterDiff = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_counterDiff : compareStage_controlPipe_translated_payload_counterDiff);
  assign compareStage_controlPipe_translated_s2mPipe_payload_twiceCompValid = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_twiceCompValid : compareStage_controlPipe_translated_payload_twiceCompValid);
  assign compareStage_controlPipe_translated_s2mPipe_payload_twiceMode = (compareStage_controlPipe_translated_rValid ? compareStage_controlPipe_translated_rData_twiceMode : compareStage_controlPipe_translated_payload_twiceMode);
  always @(*) begin
    compareStage_controlPipe_translated_s2mPipe_ready = diffStage_controlPipe_ready;
    if(when_Stream_l368_20) begin
      compareStage_controlPipe_translated_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_20 = (! diffStage_controlPipe_valid);
  assign diffStage_controlPipe_valid = compareStage_controlPipe_translated_s2mPipe_rValid;
  assign diffStage_controlPipe_payload_frameStart = compareStage_controlPipe_translated_s2mPipe_rData_frameStart;
  assign diffStage_controlPipe_payload_rowEnd = compareStage_controlPipe_translated_s2mPipe_rData_rowEnd;
  assign diffStage_controlPipe_payload_passMode = compareStage_controlPipe_translated_s2mPipe_rData_passMode;
  assign diffStage_controlPipe_payload_passValid = compareStage_controlPipe_translated_s2mPipe_rData_passValid;
  assign diffStage_controlPipe_payload_onceMode = compareStage_controlPipe_translated_s2mPipe_rData_onceMode;
  assign diffStage_controlPipe_payload_onceValid = compareStage_controlPipe_translated_s2mPipe_rData_onceValid;
  assign diffStage_controlPipe_payload_mainCompare = compareStage_controlPipe_translated_s2mPipe_rData_mainCompare;
  assign diffStage_controlPipe_payload_counterCompare = compareStage_controlPipe_translated_s2mPipe_rData_counterCompare;
  assign diffStage_controlPipe_payload_mainDiff = compareStage_controlPipe_translated_s2mPipe_rData_mainDiff;
  assign diffStage_controlPipe_payload_counterDiff = compareStage_controlPipe_translated_s2mPipe_rData_counterDiff;
  assign diffStage_controlPipe_payload_twiceCompValid = compareStage_controlPipe_translated_s2mPipe_rData_twiceCompValid;
  assign diffStage_controlPipe_payload_twiceMode = compareStage_controlPipe_translated_s2mPipe_rData_twiceMode;
  assign diffStage_mainOnePixelStream_ready = (! diffStage_mainOnePixelStream_rValid);
  assign diffStage_mainOnePixelStream_s2mPipe_valid = (diffStage_mainOnePixelStream_valid || diffStage_mainOnePixelStream_rValid);
  assign diffStage_mainOnePixelStream_s2mPipe_payload = (diffStage_mainOnePixelStream_rValid ? diffStage_mainOnePixelStream_rData : diffStage_mainOnePixelStream_payload);
  always @(*) begin
    diffStage_mainOnePixelStream_s2mPipe_ready = resultStage_mainOnePixelStream_ready;
    if(when_Stream_l368_21) begin
      diffStage_mainOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_21 = (! resultStage_mainOnePixelStream_valid);
  assign resultStage_mainOnePixelStream_valid = diffStage_mainOnePixelStream_s2mPipe_rValid;
  assign resultStage_mainOnePixelStream_payload = diffStage_mainOnePixelStream_s2mPipe_rData;
  assign diffStage_counterOnePixelStream_ready = (! diffStage_counterOnePixelStream_rValid);
  assign diffStage_counterOnePixelStream_s2mPipe_valid = (diffStage_counterOnePixelStream_valid || diffStage_counterOnePixelStream_rValid);
  assign diffStage_counterOnePixelStream_s2mPipe_payload = (diffStage_counterOnePixelStream_rValid ? diffStage_counterOnePixelStream_rData : diffStage_counterOnePixelStream_payload);
  always @(*) begin
    diffStage_counterOnePixelStream_s2mPipe_ready = resultStage_counterOnePixelStream_ready;
    if(when_Stream_l368_22) begin
      diffStage_counterOnePixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_22 = (! resultStage_counterOnePixelStream_valid);
  assign resultStage_counterOnePixelStream_valid = diffStage_counterOnePixelStream_s2mPipe_rValid;
  assign resultStage_counterOnePixelStream_payload = diffStage_counterOnePixelStream_s2mPipe_rData;
  assign diffStage_mainTwoPixelStream_ready = (! diffStage_mainTwoPixelStream_rValid);
  assign diffStage_mainTwoPixelStream_s2mPipe_valid = (diffStage_mainTwoPixelStream_valid || diffStage_mainTwoPixelStream_rValid);
  assign diffStage_mainTwoPixelStream_s2mPipe_payload = (diffStage_mainTwoPixelStream_rValid ? diffStage_mainTwoPixelStream_rData : diffStage_mainTwoPixelStream_payload);
  always @(*) begin
    diffStage_mainTwoPixelStream_s2mPipe_ready = resultStage_mainTwoPixelStream_ready;
    if(when_Stream_l368_23) begin
      diffStage_mainTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_23 = (! resultStage_mainTwoPixelStream_valid);
  assign resultStage_mainTwoPixelStream_valid = diffStage_mainTwoPixelStream_s2mPipe_rValid;
  assign resultStage_mainTwoPixelStream_payload = diffStage_mainTwoPixelStream_s2mPipe_rData;
  assign diffStage_counterTwoPixelStream_ready = (! diffStage_counterTwoPixelStream_rValid);
  assign diffStage_counterTwoPixelStream_s2mPipe_valid = (diffStage_counterTwoPixelStream_valid || diffStage_counterTwoPixelStream_rValid);
  assign diffStage_counterTwoPixelStream_s2mPipe_payload = (diffStage_counterTwoPixelStream_rValid ? diffStage_counterTwoPixelStream_rData : diffStage_counterTwoPixelStream_payload);
  always @(*) begin
    diffStage_counterTwoPixelStream_s2mPipe_ready = resultStage_counterTwoPixelStream_ready;
    if(when_Stream_l368_24) begin
      diffStage_counterTwoPixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_24 = (! resultStage_counterTwoPixelStream_valid);
  assign resultStage_counterTwoPixelStream_valid = diffStage_counterTwoPixelStream_s2mPipe_rValid;
  assign resultStage_counterTwoPixelStream_payload = diffStage_counterTwoPixelStream_s2mPipe_rData;
  assign diffStage_controlPipe_ready = diffStage_controlPipe_fork_io_input_ready;
  assign diffStage_controlPipe_fork_io_outputs_0_ready = (! diffStage_controlPipe_fork_io_outputs_0_rValid);
  assign diffStage_controlPipe_fork_io_outputs_0_s2mPipe_valid = (diffStage_controlPipe_fork_io_outputs_0_valid || diffStage_controlPipe_fork_io_outputs_0_rValid);
  assign diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_frameStart = (diffStage_controlPipe_fork_io_outputs_0_rValid ? diffStage_controlPipe_fork_io_outputs_0_rData_frameStart : diffStage_controlPipe_fork_io_outputs_0_payload_frameStart);
  assign diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_rowEnd = (diffStage_controlPipe_fork_io_outputs_0_rValid ? diffStage_controlPipe_fork_io_outputs_0_rData_rowEnd : diffStage_controlPipe_fork_io_outputs_0_payload_rowEnd);
  assign diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_passMode = (diffStage_controlPipe_fork_io_outputs_0_rValid ? diffStage_controlPipe_fork_io_outputs_0_rData_passMode : diffStage_controlPipe_fork_io_outputs_0_payload_passMode);
  assign diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_passValid = (diffStage_controlPipe_fork_io_outputs_0_rValid ? diffStage_controlPipe_fork_io_outputs_0_rData_passValid : diffStage_controlPipe_fork_io_outputs_0_payload_passValid);
  assign diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_onceMode = (diffStage_controlPipe_fork_io_outputs_0_rValid ? diffStage_controlPipe_fork_io_outputs_0_rData_onceMode : diffStage_controlPipe_fork_io_outputs_0_payload_onceMode);
  assign diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_onceValid = (diffStage_controlPipe_fork_io_outputs_0_rValid ? diffStage_controlPipe_fork_io_outputs_0_rData_onceValid : diffStage_controlPipe_fork_io_outputs_0_payload_onceValid);
  assign diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_mainCompare = (diffStage_controlPipe_fork_io_outputs_0_rValid ? diffStage_controlPipe_fork_io_outputs_0_rData_mainCompare : diffStage_controlPipe_fork_io_outputs_0_payload_mainCompare);
  assign diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_counterCompare = (diffStage_controlPipe_fork_io_outputs_0_rValid ? diffStage_controlPipe_fork_io_outputs_0_rData_counterCompare : diffStage_controlPipe_fork_io_outputs_0_payload_counterCompare);
  assign diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_mainDiff = (diffStage_controlPipe_fork_io_outputs_0_rValid ? diffStage_controlPipe_fork_io_outputs_0_rData_mainDiff : diffStage_controlPipe_fork_io_outputs_0_payload_mainDiff);
  assign diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_counterDiff = (diffStage_controlPipe_fork_io_outputs_0_rValid ? diffStage_controlPipe_fork_io_outputs_0_rData_counterDiff : diffStage_controlPipe_fork_io_outputs_0_payload_counterDiff);
  assign diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_twiceCompValid = (diffStage_controlPipe_fork_io_outputs_0_rValid ? diffStage_controlPipe_fork_io_outputs_0_rData_twiceCompValid : diffStage_controlPipe_fork_io_outputs_0_payload_twiceCompValid);
  assign diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_twiceMode = (diffStage_controlPipe_fork_io_outputs_0_rValid ? diffStage_controlPipe_fork_io_outputs_0_rData_twiceMode : diffStage_controlPipe_fork_io_outputs_0_payload_twiceMode);
  always @(*) begin
    diffStage_controlPipe_fork_io_outputs_0_s2mPipe_ready = resultStage_controlPipe_ready;
    if(when_Stream_l368_25) begin
      diffStage_controlPipe_fork_io_outputs_0_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_25 = (! resultStage_controlPipe_valid);
  assign resultStage_controlPipe_valid = diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rValid;
  assign resultStage_controlPipe_payload_frameStart = diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_frameStart;
  assign resultStage_controlPipe_payload_rowEnd = diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_rowEnd;
  assign resultStage_controlPipe_payload_passMode = diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_passMode;
  assign resultStage_controlPipe_payload_passValid = diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_passValid;
  assign resultStage_controlPipe_payload_onceMode = diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_onceMode;
  assign resultStage_controlPipe_payload_onceValid = diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_onceValid;
  assign resultStage_controlPipe_payload_mainCompare = diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_mainCompare;
  assign resultStage_controlPipe_payload_counterCompare = diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_counterCompare;
  assign resultStage_controlPipe_payload_mainDiff = diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_mainDiff;
  assign resultStage_controlPipe_payload_counterDiff = diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_counterDiff;
  assign resultStage_controlPipe_payload_twiceCompValid = diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_twiceCompValid;
  assign resultStage_controlPipe_payload_twiceMode = diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_twiceMode;
  assign resultStage_pixelStream_valid = diffStage_controlPipe_fork_io_outputs_1_valid;
  always @(*) begin
    resultStage_pixelStream_payload = 8'h0;
    if(diffStage_controlPipe_fork_io_outputs_1_payload_passValid) begin
      if(diffStage_controlPipe_fork_io_outputs_1_payload_passMode) begin
        resultStage_pixelStream_payload = diffStage_mainTwoPixelStream_payload;
      end else begin
        resultStage_pixelStream_payload = diffStage_mainOnePixelStream_payload;
      end
    end
    if(diffStage_controlPipe_fork_io_outputs_1_payload_onceValid) begin
      case(diffStage_controlPipe_fork_io_outputs_1_payload_onceMode)
        3'b000 : begin
          if(when_SuperResolutionPart1_l339) begin
            resultStage_pixelStream_payload = diffStage_mainOnePixelStream_payload;
          end else begin
            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload[7:0];
          end
        end
        3'b001 : begin
          if(when_SuperResolutionPart1_l343) begin
            resultStage_pixelStream_payload = diffStage_mainTwoPixelStream_payload;
          end else begin
            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_2[7:0];
          end
        end
        3'b010 : begin
          if(when_SuperResolutionPart1_l347) begin
            resultStage_pixelStream_payload = diffStage_mainOnePixelStream_payload;
          end else begin
            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_4[7:0];
          end
        end
        3'b011 : begin
          if(when_SuperResolutionPart1_l351) begin
            resultStage_pixelStream_payload = diffStage_mainTwoPixelStream_payload;
          end else begin
            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_6[7:0];
          end
        end
        3'b100 : begin
          resultStage_pixelStream_payload = diffStage_mainTwoPixelStream_payload;
        end
        3'b101 : begin
          resultStage_pixelStream_payload = diffStage_mainOnePixelStream_payload;
        end
        default : begin
        end
      endcase
    end
    if(diffStage_controlPipe_fork_io_outputs_1_payload_twiceCompValid) begin
      case(diffStage_controlPipe_fork_io_outputs_1_payload_twiceMode)
        3'b000 : begin
          if(when_SuperResolutionPart1_l362) begin
            if(when_SuperResolutionPart1_l363) begin
              resultStage_pixelStream_payload = diffStage_mainOnePixelStream_payload;
            end else begin
              resultStage_pixelStream_payload = diffStage_counterTwoPixelStream_payload;
            end
          end else begin
            if(when_SuperResolutionPart1_l366) begin
              resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_8[7:0];
            end else begin
              resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_10[7:0];
            end
          end
        end
        3'b001 : begin
          if(when_SuperResolutionPart1_l371) begin
            if(when_SuperResolutionPart1_l372) begin
              resultStage_pixelStream_payload = diffStage_mainTwoPixelStream_payload;
            end else begin
              resultStage_pixelStream_payload = diffStage_counterOnePixelStream_payload;
            end
          end else begin
            if(when_SuperResolutionPart1_l375) begin
              resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_12[7:0];
            end else begin
              resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_14[7:0];
            end
          end
        end
        3'b010 : begin
          resultStage_pixelStream_payload = diffStage_mainTwoPixelStream_payload;
        end
        3'b011 : begin
          if(when_SuperResolutionPart1_l381) begin
            resultStage_pixelStream_payload = diffStage_mainTwoPixelStream_payload;
          end else begin
            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_16[7:0];
          end
        end
        3'b100 : begin
          resultStage_pixelStream_payload = diffStage_mainOnePixelStream_payload;
        end
        3'b101 : begin
          if(when_SuperResolutionPart1_l386) begin
            resultStage_pixelStream_payload = diffStage_mainOnePixelStream_payload;
          end else begin
            resultStage_pixelStream_payload = CICC1851_resultStage_pixelStream_payload_18[7:0];
          end
        end
        default : begin
        end
      endcase
    end
  end

  assign when_SuperResolutionPart1_l339 = (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart1_l343 = (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart1_l347 = (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart1_l351 = (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart1_l362 = ((inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff) && (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff));
  assign when_SuperResolutionPart1_l363 = (diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart1_l366 = (diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart1_l371 = ((inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff) && (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff));
  assign when_SuperResolutionPart1_l372 = (diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart1_l375 = (diffStage_controlPipe_fork_io_outputs_1_payload_counterDiff <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart1_l381 = (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign when_SuperResolutionPart1_l386 = (inpThreshold <= diffStage_controlPipe_fork_io_outputs_1_payload_mainDiff);
  assign resultStage_pixelStream_ready = (! resultStage_pixelStream_rValid);
  assign resultStage_pixelStream_s2mPipe_valid = (resultStage_pixelStream_valid || resultStage_pixelStream_rValid);
  assign resultStage_pixelStream_s2mPipe_payload = (resultStage_pixelStream_rValid ? resultStage_pixelStream_rData : resultStage_pixelStream_payload);
  always @(*) begin
    resultStage_pixelStream_s2mPipe_ready = resultStage_resultStream_ready;
    if(when_Stream_l368_26) begin
      resultStage_pixelStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_26 = (! resultStage_resultStream_valid);
  assign resultStage_resultStream_valid = resultStage_pixelStream_s2mPipe_rValid;
  assign resultStage_resultStream_payload = resultStage_pixelStream_s2mPipe_rData;
  assign CICC1851_resultStage_mainOnePixelStream_ready_2 = (CICC1851_resultStage_mainOnePixelStream_ready && CICC1851_resultStage_mainOnePixelStream_ready_1);
  assign CICC1851_resultStage_mainOnePixelStream_ready = (((((resultStage_resultStream_valid && resultStage_mainOnePixelStream_valid) && resultStage_counterOnePixelStream_valid) && resultStage_mainTwoPixelStream_valid) && resultStage_counterTwoPixelStream_valid) && resultStage_controlPipe_valid);
  assign resultStage_resultStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_mainOnePixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_counterOnePixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_mainTwoPixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_counterTwoPixelStream_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign resultStage_controlPipe_ready = CICC1851_resultStage_mainOnePixelStream_ready_2;
  assign when_Stream_l438 = (((! resultStage_controlPipe_payload_passValid) && (! resultStage_controlPipe_payload_onceValid)) && (! resultStage_controlPipe_payload_twiceCompValid));
  always @(*) begin
    resultsJoin_valid = CICC1851_resultStage_mainOnePixelStream_ready;
    if(when_Stream_l438) begin
      resultsJoin_valid = 1'b0;
    end
  end

  always @(*) begin
    CICC1851_resultStage_mainOnePixelStream_ready_1 = resultsJoin_ready;
    if(when_Stream_l438) begin
      CICC1851_resultStage_mainOnePixelStream_ready_1 = 1'b1;
    end
  end

  assign pixelsStream_valid = resultsJoin_valid;
  assign resultsJoin_ready = pixelsStream_ready;
  assign pixelsStream_payload_pixel = resultStage_resultStream_payload;
  assign pixelsStream_payload_frameStart = resultStage_controlPipe_payload_frameStart;
  assign pixelsStream_payload_rowEnd = resultStage_controlPipe_payload_rowEnd;
  assign pixelsStream_ready = (! pixelsStream_rValid);
  assign pixelsStream_s2mPipe_valid = (pixelsStream_valid || pixelsStream_rValid);
  assign pixelsStream_s2mPipe_payload_pixel = (pixelsStream_rValid ? pixelsStream_rData_pixel : pixelsStream_payload_pixel);
  assign pixelsStream_s2mPipe_payload_frameStart = (pixelsStream_rValid ? pixelsStream_rData_frameStart : pixelsStream_payload_frameStart);
  assign pixelsStream_s2mPipe_payload_rowEnd = (pixelsStream_rValid ? pixelsStream_rData_rowEnd : pixelsStream_payload_rowEnd);
  always @(*) begin
    pixelsStream_s2mPipe_ready = pixelsStream_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_27) begin
      pixelsStream_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_27 = (! pixelsStream_s2mPipe_m2sPipe_valid);
  assign pixelsStream_s2mPipe_m2sPipe_valid = pixelsStream_s2mPipe_rValid;
  assign pixelsStream_s2mPipe_m2sPipe_payload_pixel = pixelsStream_s2mPipe_rData_pixel;
  assign pixelsStream_s2mPipe_m2sPipe_payload_frameStart = pixelsStream_s2mPipe_rData_frameStart;
  assign pixelsStream_s2mPipe_m2sPipe_payload_rowEnd = pixelsStream_s2mPipe_rData_rowEnd;
  assign pixelsStream_s2mPipe_m2sPipe_ready = pixelsOut_ready;
  assign pixelsIn_s2mPipe_valid = (pixelsIn_valid || pixelsIn_rValid);
  assign pixelsIn_s2mPipe_payload_pixel = (pixelsIn_rValid ? pixelsIn_rData_pixel : pixelsIn_payload_pixel);
  assign pixelsIn_s2mPipe_payload_frameStart = (pixelsIn_rValid ? pixelsIn_rData_frameStart : pixelsIn_payload_frameStart);
  assign pixelsIn_s2mPipe_payload_rowEnd = (pixelsIn_rValid ? pixelsIn_rData_rowEnd : pixelsIn_payload_rowEnd);
  always @(*) begin
    pixelsIn_s2mPipe_ready = pixelsIn_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_28) begin
      pixelsIn_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_28 = (! pixelsIn_s2mPipe_m2sPipe_valid);
  assign pixelsIn_s2mPipe_m2sPipe_valid = pixelsIn_s2mPipe_rValid;
  assign pixelsIn_s2mPipe_m2sPipe_payload_pixel = pixelsIn_s2mPipe_rData_pixel;
  assign pixelsIn_s2mPipe_m2sPipe_payload_frameStart = pixelsIn_s2mPipe_rData_frameStart;
  assign pixelsIn_s2mPipe_m2sPipe_payload_rowEnd = pixelsIn_s2mPipe_rData_rowEnd;
  assign passPixels_valid = (pixelsIn_s2mPipe_m2sPipe_valid && bufferEnable);
  assign pixelsIn_s2mPipe_m2sPipe_ready = (passPixels_ready && bufferEnable);
  assign passPixels_payload_pixel = pixelsIn_s2mPipe_m2sPipe_payload_pixel;
  assign passPixels_payload_frameStart = pixelsIn_s2mPipe_m2sPipe_payload_frameStart;
  assign passPixels_payload_rowEnd = pixelsIn_s2mPipe_m2sPipe_payload_rowEnd;
  assign passPixels_ready = 1'b1;
  assign passPixels_fire = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart1_l421 = ((bufferWAddr_value == CICC1851_when_SuperResolutionPart1_l421) && passPixels_fire);
  assign passPixels_fire_1 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart1_l422 = (((bufferRowCount_value == CICC1851_when_SuperResolutionPart1_l422) && bufferReachRowEnd) && passPixels_fire_1);
  assign passPixels_fire_2 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart1_l425 = (passPixels_payload_rowEnd && passPixels_fire_2);
  assign passPixels_fire_3 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart1_l438 = (passPixels_payload_rowEnd && passPixels_fire_3);
  assign passPixels_fire_4 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart1_l439 = (((bufferRowCount_value != 10'h0) && passPixels_payload_rowEnd) && passPixels_fire_4);
  assign when_SuperResolutionPart1_l442 = (bufferReachFinalRow && bufferReachRowEnd);
  assign controlStream_fire = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l447 = (((CICC1851_when_SuperResolutionPart1_l447 == 11'h001) && controlStream_payload_rowEnd) && controlStream_fire);
  assign when_SuperResolutionPart1_l449 = 1'b1;
  assign passPixels_fire_5 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart1_l453 = (passPixels_payload_frameStart && passPixels_fire_5);
  assign passPixels_fire_6 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_7 = (passPixels_valid && passPixels_ready);
  assign passPixels_fire_8 = (passPixels_valid && passPixels_ready);
  assign controlStateMachine_wantExit = 1'b0;
  always @(*) begin
    controlStateMachine_wantStart = 1'b0;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_HOLD : begin
      end
      controlStateMachine_enumDef_PASS : begin
      end
      controlStateMachine_enumDef_ONCE : begin
      end
      controlStateMachine_enumDef_TWICE : begin
      end
      default : begin
        controlStateMachine_wantStart = 1'b1;
      end
    endcase
  end

  assign controlStateMachine_wantKill = 1'b0;
  always @(*) begin
    controlStateMachine_stateNext = controlStateMachine_stateReg;
    case(controlStateMachine_stateReg)
      controlStateMachine_enumDef_HOLD : begin
        if(when_SuperResolutionPart1_l482) begin
          if(passPixels_fire_9) begin
            if(when_SuperResolutionPart1_l484) begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_PASS;
            end else begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_ONCE;
            end
          end
        end else begin
          if(passPixels_fire_10) begin
            if(when_SuperResolutionPart1_l489) begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_ONCE;
            end else begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_TWICE;
            end
          end
        end
      end
      controlStateMachine_enumDef_PASS : begin
        if(controlStream_fire_1) begin
          if(when_SuperResolutionPart1_l498) begin
            controlStateMachine_stateNext = controlStateMachine_enumDef_ONCE;
          end else begin
            if(when_SuperResolutionPart1_l500) begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_HOLD;
            end else begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_ONCE;
            end
          end
        end
      end
      controlStateMachine_enumDef_ONCE : begin
        if(when_SuperResolutionPart1_l537) begin
          if(controlStream_fire_7) begin
            if(outReachRowEnd) begin
              if(bufferReuse) begin
                controlStateMachine_stateNext = controlStateMachine_enumDef_ONCE;
              end else begin
                if(when_SuperResolutionPart1_l542) begin
                  controlStateMachine_stateNext = controlStateMachine_enumDef_HOLD;
                end else begin
                  controlStateMachine_stateNext = controlStateMachine_enumDef_ONCE;
                end
              end
            end else begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_PASS;
            end
          end
        end else begin
          if(controlStream_fire_8) begin
            if(bufferReuse) begin
              controlStateMachine_stateNext = controlStateMachine_enumDef_TWICE;
            end else begin
              if(when_SuperResolutionPart1_l563) begin
                controlStateMachine_stateNext = controlStateMachine_enumDef_HOLD;
              end else begin
                controlStateMachine_stateNext = controlStateMachine_enumDef_TWICE;
              end
            end
          end
        end
      end
      controlStateMachine_enumDef_TWICE : begin
        if(controlStream_fire_13) begin
          if(outReachRowEnd) begin
            if(bufferReuse) begin
              if(outReachFinalRow) begin
                controlStateMachine_stateNext = controlStateMachine_enumDef_HOLD;
              end else begin
                controlStateMachine_stateNext = controlStateMachine_enumDef_PASS;
              end
            end else begin
              if(when_SuperResolutionPart1_l612) begin
                controlStateMachine_stateNext = controlStateMachine_enumDef_HOLD;
              end else begin
                controlStateMachine_stateNext = controlStateMachine_enumDef_PASS;
              end
            end
          end else begin
            controlStateMachine_stateNext = controlStateMachine_enumDef_ONCE;
          end
        end
      end
      default : begin
      end
    endcase
    if(controlStateMachine_wantStart) begin
      controlStateMachine_stateNext = controlStateMachine_enumDef_HOLD;
    end
    if(controlStateMachine_wantKill) begin
      controlStateMachine_stateNext = controlStateMachine_enumDef_BOOT;
    end
  end

  assign when_SuperResolutionPart1_l482 = (CICC1851_when_SuperResolutionPart1_l482 == 11'h0);
  assign passPixels_fire_9 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart1_l484 = (CICC1851_when_SuperResolutionPart1_l484 == 11'h0);
  assign passPixels_fire_10 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart1_l489 = (CICC1851_when_SuperResolutionPart1_l489 == 11'h0);
  assign controlStream_fire_1 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l498 = ((CICC1851_when_SuperResolutionPart1_l498 < CICC1851_when_SuperResolutionPart1_l498_1) || bufferReuse);
  assign passPixels_fire_11 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart1_l500 = ((CICC1851_when_SuperResolutionPart1_l500 == CICC1851_when_SuperResolutionPart1_l500_1) && (! passPixels_fire_11));
  assign controlStream_fire_2 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l507 = (frameStart && controlStream_fire_2);
  assign controlStream_fire_3 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l510 = (controlStream_fire_3 && (CICC1851_when_SuperResolutionPart1_l510 == CICC1851_when_SuperResolutionPart1_l510_1));
  assign controlStream_fire_4 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l511 = ((outReachRowEnd && (CICC1851_when_SuperResolutionPart1_l511 == CICC1851_when_SuperResolutionPart1_l511_1)) && controlStream_fire_4);
  assign controlStream_fire_5 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l513 = (controlStream_fire_5 && outReachRowEnd);
  assign controlStream_fire_6 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l537 = (CICC1851_when_SuperResolutionPart1_l537 == 11'h0);
  assign controlStream_fire_7 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l542 = ((bufferWAddr_value == 10'h0) && (CICC1851_when_SuperResolutionPart1_l542 == CICC1851_when_SuperResolutionPart1_l542_2));
  assign controlStream_fire_8 = (controlStream_valid && controlStream_ready);
  assign passPixels_fire_12 = (passPixels_valid && passPixels_ready);
  assign when_SuperResolutionPart1_l563 = ((CICC1851_when_SuperResolutionPart1_l563 == CICC1851_when_SuperResolutionPart1_l563_1) && (! passPixels_fire_12));
  assign controlStream_fire_9 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l578 = (controlStream_fire_9 && (CICC1851_when_SuperResolutionPart1_l578 == CICC1851_when_SuperResolutionPart1_l578_1));
  assign controlStream_fire_10 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l579 = ((outReachRowEnd && (CICC1851_when_SuperResolutionPart1_l579 == CICC1851_when_SuperResolutionPart1_l579_1)) && controlStream_fire_10);
  assign controlStream_fire_11 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l581 = (controlStream_fire_11 && outReachRowEnd);
  assign controlStream_fire_12 = (controlStream_valid && controlStream_ready);
  assign controlStream_fire_13 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l612 = (bufferWAddr_value == 10'h0);
  assign controlStream_fire_14 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l664 = (controlStream_fire_14 && (CICC1851_when_SuperResolutionPart1_l664 == CICC1851_when_SuperResolutionPart1_l664_1));
  assign controlStream_fire_15 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l665 = ((outReachRowEnd && (CICC1851_when_SuperResolutionPart1_l665 == CICC1851_when_SuperResolutionPart1_l665_1)) && controlStream_fire_15);
  assign controlStream_fire_16 = (controlStream_valid && controlStream_ready);
  assign when_SuperResolutionPart1_l667 = (controlStream_fire_16 && outReachRowEnd);
  assign controlStream_fire_17 = (controlStream_valid && controlStream_ready);
  always @(posedge clk or negedge resetn) begin
    if(!resetn) begin
      inpDone <= 1'b0;
      readDone <= 1'b0;
      startRead <= 1'b0;
      slaveStart <= 1'b0;
      frameStart <= 1'b0;
      inpThreshold <= 8'h80;
      bmpWidth <= 10'h3c0;
      bmpHeight <= 10'h21c;
      holdBuffer <= 1'b0;
      writeDone <= 1'b0;
      bufferRowCount_value <= 10'h0;
      bufferEnable <= 1'b0;
      bufferSwitch <= 1'b0;
      nextRowBuffer <= 1'b1;
      bufferReuse <= 1'b0;
      bufferWAddr_value <= 10'h0;
      outPixelAddr_value <= 11'h0;
      outRowCount_value <= 11'h0;
      outReachRowEnd <= 1'b0;
      outReachFinalRow <= 1'b0;
      bufferReachRowEnd <= 1'b0;
      bufferReachFinalRow <= 1'b0;
      mainAddrOneStream_rValid <= 1'b0;
      mainAddrOneStream_s2mPipe_rValid <= 1'b0;
      CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_mainOnePixelStream_valid <= 1'b0;
      counterAddrOneStream_rValid <= 1'b0;
      counterAddrOneStream_s2mPipe_rValid <= 1'b0;
      CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_counterOnePixelStream_valid <= 1'b0;
      mainAddrTwoStream_rValid <= 1'b0;
      mainAddrTwoStream_s2mPipe_rValid <= 1'b0;
      CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_mainTwoPixelStream_valid <= 1'b0;
      counterAddrTwoStream_rValid <= 1'b0;
      counterAddrTwoStream_s2mPipe_rValid <= 1'b0;
      CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      CICC1851_readStage_counterTwoPixelStream_valid <= 1'b0;
      controlStream_rValid <= 1'b0;
      controlStream_s2mPipe_rValid <= 1'b0;
      controlStream_s2mPipe_m2sPipe_rValid <= 1'b0;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rValid <= 1'b0;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rValid <= 1'b0;
      readStage_mainOnePixelStream_rValid <= 1'b0;
      readStage_mainOnePixelStream_s2mPipe_rValid <= 1'b0;
      readStage_counterOnePixelStream_rValid <= 1'b0;
      readStage_counterOnePixelStream_s2mPipe_rValid <= 1'b0;
      readStage_mainTwoPixelStream_rValid <= 1'b0;
      readStage_mainTwoPixelStream_s2mPipe_rValid <= 1'b0;
      readStage_counterTwoPixelStream_rValid <= 1'b0;
      readStage_counterTwoPixelStream_s2mPipe_rValid <= 1'b0;
      readStage_controlPipe_translated_rValid <= 1'b0;
      readStage_controlPipe_translated_s2mPipe_rValid <= 1'b0;
      compareStage_mainOnePixelStream_rValid <= 1'b0;
      compareStage_mainOnePixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_counterOnePixelStream_rValid <= 1'b0;
      compareStage_counterOnePixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_mainTwoPixelStream_rValid <= 1'b0;
      compareStage_mainTwoPixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_counterTwoPixelStream_rValid <= 1'b0;
      compareStage_counterTwoPixelStream_s2mPipe_rValid <= 1'b0;
      compareStage_controlPipe_translated_rValid <= 1'b0;
      compareStage_controlPipe_translated_s2mPipe_rValid <= 1'b0;
      diffStage_mainOnePixelStream_rValid <= 1'b0;
      diffStage_mainOnePixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_counterOnePixelStream_rValid <= 1'b0;
      diffStage_counterOnePixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_mainTwoPixelStream_rValid <= 1'b0;
      diffStage_mainTwoPixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_counterTwoPixelStream_rValid <= 1'b0;
      diffStage_counterTwoPixelStream_s2mPipe_rValid <= 1'b0;
      diffStage_controlPipe_fork_io_outputs_0_rValid <= 1'b0;
      diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rValid <= 1'b0;
      resultStage_pixelStream_rValid <= 1'b0;
      resultStage_pixelStream_s2mPipe_rValid <= 1'b0;
      pixelsStream_rValid <= 1'b0;
      pixelsStream_s2mPipe_rValid <= 1'b0;
      pixelsIn_rValid <= 1'b0;
      pixelsIn_s2mPipe_rValid <= 1'b0;
      controlStateMachine_stateReg <= controlStateMachine_enumDef_BOOT;
    end else begin
      if(when_SuperResolutionPart1_l79) begin
        inpDone <= 1'b1;
      end
      if(when_SuperResolutionPart1_l79_1) begin
        inpDone <= 1'b0;
      end
      if(when_SuperResolutionPart1_l82) begin
        readDone <= 1'b0;
      end
      if(when_SuperResolutionPart1_l85) begin
        startRead <= 1'b1;
      end
      if(when_SuperResolutionPart1_l85_1) begin
        startRead <= 1'b0;
      end
      if(when_SuperResolutionPart1_l88) begin
        slaveStart <= 1'b1;
      end
      if(when_SuperResolutionPart1_l88_1) begin
        slaveStart <= 1'b0;
      end
      inpThreshold <= thresholdIn;
      bmpWidth <= widthIn;
      bmpHeight <= heightIn;
      if(when_SuperResolutionPart1_l103) begin
        holdBuffer <= 1'b0;
      end
      if(when_SuperResolutionPart1_l106) begin
        writeDone <= 1'b0;
      end
      bufferRowCount_value <= bufferRowCount_valueNext;
      if(when_SuperResolutionPart1_l112) begin
        bufferEnable <= 1'b1;
      end
      if(when_SuperResolutionPart1_l112_1) begin
        bufferEnable <= 1'b0;
      end
      if(when_SuperResolutionPart1_l115) begin
        bufferSwitch <= 1'b0;
      end
      if(when_SuperResolutionPart1_l118) begin
        nextRowBuffer <= 1'b1;
      end
      if(inpDone) begin
        bufferReuse <= 1'b0;
      end
      bufferWAddr_value <= bufferWAddr_valueNext;
      outPixelAddr_value <= outPixelAddr_valueNext;
      outRowCount_value <= outRowCount_valueNext;
      if(mainAddrOneStream_valid) begin
        mainAddrOneStream_rValid <= 1'b1;
      end
      if(mainAddrOneStream_s2mPipe_ready) begin
        mainAddrOneStream_rValid <= 1'b0;
      end
      if(mainAddrOneStream_s2mPipe_ready) begin
        mainAddrOneStream_s2mPipe_rValid <= mainAddrOneStream_s2mPipe_valid;
      end
      if(CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(mainAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_2 <= mainAddrOneStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_1) begin
        CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_1) begin
        CICC1851_readStage_mainOnePixelStream_valid <= (CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready || CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_3);
      end
      if(counterAddrOneStream_valid) begin
        counterAddrOneStream_rValid <= 1'b1;
      end
      if(counterAddrOneStream_s2mPipe_ready) begin
        counterAddrOneStream_rValid <= 1'b0;
      end
      if(counterAddrOneStream_s2mPipe_ready) begin
        counterAddrOneStream_s2mPipe_rValid <= counterAddrOneStream_s2mPipe_valid;
      end
      if(CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(counterAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_2 <= counterAddrOneStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_2) begin
        CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_2) begin
        CICC1851_readStage_counterOnePixelStream_valid <= (CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready || CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_3);
      end
      if(mainAddrTwoStream_valid) begin
        mainAddrTwoStream_rValid <= 1'b1;
      end
      if(mainAddrTwoStream_s2mPipe_ready) begin
        mainAddrTwoStream_rValid <= 1'b0;
      end
      if(mainAddrTwoStream_s2mPipe_ready) begin
        mainAddrTwoStream_s2mPipe_rValid <= mainAddrTwoStream_s2mPipe_valid;
      end
      if(CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(mainAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= mainAddrTwoStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_3) begin
        CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_3) begin
        CICC1851_readStage_mainTwoPixelStream_valid <= (CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready || CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_3);
      end
      if(counterAddrTwoStream_valid) begin
        counterAddrTwoStream_rValid <= 1'b1;
      end
      if(counterAddrTwoStream_s2mPipe_ready) begin
        counterAddrTwoStream_rValid <= 1'b0;
      end
      if(counterAddrTwoStream_s2mPipe_ready) begin
        counterAddrTwoStream_s2mPipe_rValid <= counterAddrTwoStream_s2mPipe_valid;
      end
      if(CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
        CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= 1'b0;
      end
      if(counterAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_2 <= counterAddrTwoStream_s2mPipe_m2sPipe_valid;
      end
      if(CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready) begin
        CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b1;
      end
      if(CICC1851_4) begin
        CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_3 <= 1'b0;
      end
      if(CICC1851_4) begin
        CICC1851_readStage_counterTwoPixelStream_valid <= (CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready || CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_3);
      end
      if(controlStream_valid) begin
        controlStream_rValid <= 1'b1;
      end
      if(controlStream_s2mPipe_ready) begin
        controlStream_rValid <= 1'b0;
      end
      if(controlStream_s2mPipe_ready) begin
        controlStream_s2mPipe_rValid <= controlStream_s2mPipe_valid;
      end
      if(controlStream_s2mPipe_m2sPipe_ready) begin
        controlStream_s2mPipe_m2sPipe_rValid <= controlStream_s2mPipe_m2sPipe_valid;
      end
      if(controlStream_s2mPipe_m2sPipe_m2sPipe_valid) begin
        controlStream_s2mPipe_m2sPipe_m2sPipe_rValid <= 1'b1;
      end
      if(controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready) begin
        controlStream_s2mPipe_m2sPipe_m2sPipe_rValid <= 1'b0;
      end
      if(controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready) begin
        controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_valid;
      end
      if(readStage_mainOnePixelStream_valid) begin
        readStage_mainOnePixelStream_rValid <= 1'b1;
      end
      if(readStage_mainOnePixelStream_s2mPipe_ready) begin
        readStage_mainOnePixelStream_rValid <= 1'b0;
      end
      if(readStage_mainOnePixelStream_s2mPipe_ready) begin
        readStage_mainOnePixelStream_s2mPipe_rValid <= readStage_mainOnePixelStream_s2mPipe_valid;
      end
      if(readStage_counterOnePixelStream_valid) begin
        readStage_counterOnePixelStream_rValid <= 1'b1;
      end
      if(readStage_counterOnePixelStream_s2mPipe_ready) begin
        readStage_counterOnePixelStream_rValid <= 1'b0;
      end
      if(readStage_counterOnePixelStream_s2mPipe_ready) begin
        readStage_counterOnePixelStream_s2mPipe_rValid <= readStage_counterOnePixelStream_s2mPipe_valid;
      end
      if(readStage_mainTwoPixelStream_valid) begin
        readStage_mainTwoPixelStream_rValid <= 1'b1;
      end
      if(readStage_mainTwoPixelStream_s2mPipe_ready) begin
        readStage_mainTwoPixelStream_rValid <= 1'b0;
      end
      if(readStage_mainTwoPixelStream_s2mPipe_ready) begin
        readStage_mainTwoPixelStream_s2mPipe_rValid <= readStage_mainTwoPixelStream_s2mPipe_valid;
      end
      if(readStage_counterTwoPixelStream_valid) begin
        readStage_counterTwoPixelStream_rValid <= 1'b1;
      end
      if(readStage_counterTwoPixelStream_s2mPipe_ready) begin
        readStage_counterTwoPixelStream_rValid <= 1'b0;
      end
      if(readStage_counterTwoPixelStream_s2mPipe_ready) begin
        readStage_counterTwoPixelStream_s2mPipe_rValid <= readStage_counterTwoPixelStream_s2mPipe_valid;
      end
      if(readStage_controlPipe_translated_valid) begin
        readStage_controlPipe_translated_rValid <= 1'b1;
      end
      if(readStage_controlPipe_translated_s2mPipe_ready) begin
        readStage_controlPipe_translated_rValid <= 1'b0;
      end
      if(readStage_controlPipe_translated_s2mPipe_ready) begin
        readStage_controlPipe_translated_s2mPipe_rValid <= readStage_controlPipe_translated_s2mPipe_valid;
      end
      if(compareStage_mainOnePixelStream_valid) begin
        compareStage_mainOnePixelStream_rValid <= 1'b1;
      end
      if(compareStage_mainOnePixelStream_s2mPipe_ready) begin
        compareStage_mainOnePixelStream_rValid <= 1'b0;
      end
      if(compareStage_mainOnePixelStream_s2mPipe_ready) begin
        compareStage_mainOnePixelStream_s2mPipe_rValid <= compareStage_mainOnePixelStream_s2mPipe_valid;
      end
      if(compareStage_counterOnePixelStream_valid) begin
        compareStage_counterOnePixelStream_rValid <= 1'b1;
      end
      if(compareStage_counterOnePixelStream_s2mPipe_ready) begin
        compareStage_counterOnePixelStream_rValid <= 1'b0;
      end
      if(compareStage_counterOnePixelStream_s2mPipe_ready) begin
        compareStage_counterOnePixelStream_s2mPipe_rValid <= compareStage_counterOnePixelStream_s2mPipe_valid;
      end
      if(compareStage_mainTwoPixelStream_valid) begin
        compareStage_mainTwoPixelStream_rValid <= 1'b1;
      end
      if(compareStage_mainTwoPixelStream_s2mPipe_ready) begin
        compareStage_mainTwoPixelStream_rValid <= 1'b0;
      end
      if(compareStage_mainTwoPixelStream_s2mPipe_ready) begin
        compareStage_mainTwoPixelStream_s2mPipe_rValid <= compareStage_mainTwoPixelStream_s2mPipe_valid;
      end
      if(compareStage_counterTwoPixelStream_valid) begin
        compareStage_counterTwoPixelStream_rValid <= 1'b1;
      end
      if(compareStage_counterTwoPixelStream_s2mPipe_ready) begin
        compareStage_counterTwoPixelStream_rValid <= 1'b0;
      end
      if(compareStage_counterTwoPixelStream_s2mPipe_ready) begin
        compareStage_counterTwoPixelStream_s2mPipe_rValid <= compareStage_counterTwoPixelStream_s2mPipe_valid;
      end
      if(compareStage_controlPipe_translated_valid) begin
        compareStage_controlPipe_translated_rValid <= 1'b1;
      end
      if(compareStage_controlPipe_translated_s2mPipe_ready) begin
        compareStage_controlPipe_translated_rValid <= 1'b0;
      end
      if(compareStage_controlPipe_translated_s2mPipe_ready) begin
        compareStage_controlPipe_translated_s2mPipe_rValid <= compareStage_controlPipe_translated_s2mPipe_valid;
      end
      if(diffStage_mainOnePixelStream_valid) begin
        diffStage_mainOnePixelStream_rValid <= 1'b1;
      end
      if(diffStage_mainOnePixelStream_s2mPipe_ready) begin
        diffStage_mainOnePixelStream_rValid <= 1'b0;
      end
      if(diffStage_mainOnePixelStream_s2mPipe_ready) begin
        diffStage_mainOnePixelStream_s2mPipe_rValid <= diffStage_mainOnePixelStream_s2mPipe_valid;
      end
      if(diffStage_counterOnePixelStream_valid) begin
        diffStage_counterOnePixelStream_rValid <= 1'b1;
      end
      if(diffStage_counterOnePixelStream_s2mPipe_ready) begin
        diffStage_counterOnePixelStream_rValid <= 1'b0;
      end
      if(diffStage_counterOnePixelStream_s2mPipe_ready) begin
        diffStage_counterOnePixelStream_s2mPipe_rValid <= diffStage_counterOnePixelStream_s2mPipe_valid;
      end
      if(diffStage_mainTwoPixelStream_valid) begin
        diffStage_mainTwoPixelStream_rValid <= 1'b1;
      end
      if(diffStage_mainTwoPixelStream_s2mPipe_ready) begin
        diffStage_mainTwoPixelStream_rValid <= 1'b0;
      end
      if(diffStage_mainTwoPixelStream_s2mPipe_ready) begin
        diffStage_mainTwoPixelStream_s2mPipe_rValid <= diffStage_mainTwoPixelStream_s2mPipe_valid;
      end
      if(diffStage_counterTwoPixelStream_valid) begin
        diffStage_counterTwoPixelStream_rValid <= 1'b1;
      end
      if(diffStage_counterTwoPixelStream_s2mPipe_ready) begin
        diffStage_counterTwoPixelStream_rValid <= 1'b0;
      end
      if(diffStage_counterTwoPixelStream_s2mPipe_ready) begin
        diffStage_counterTwoPixelStream_s2mPipe_rValid <= diffStage_counterTwoPixelStream_s2mPipe_valid;
      end
      if(diffStage_controlPipe_fork_io_outputs_0_valid) begin
        diffStage_controlPipe_fork_io_outputs_0_rValid <= 1'b1;
      end
      if(diffStage_controlPipe_fork_io_outputs_0_s2mPipe_ready) begin
        diffStage_controlPipe_fork_io_outputs_0_rValid <= 1'b0;
      end
      if(diffStage_controlPipe_fork_io_outputs_0_s2mPipe_ready) begin
        diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rValid <= diffStage_controlPipe_fork_io_outputs_0_s2mPipe_valid;
      end
      if(resultStage_pixelStream_valid) begin
        resultStage_pixelStream_rValid <= 1'b1;
      end
      if(resultStage_pixelStream_s2mPipe_ready) begin
        resultStage_pixelStream_rValid <= 1'b0;
      end
      if(resultStage_pixelStream_s2mPipe_ready) begin
        resultStage_pixelStream_s2mPipe_rValid <= resultStage_pixelStream_s2mPipe_valid;
      end
      if(pixelsStream_valid) begin
        pixelsStream_rValid <= 1'b1;
      end
      if(pixelsStream_s2mPipe_ready) begin
        pixelsStream_rValid <= 1'b0;
      end
      if(pixelsStream_s2mPipe_ready) begin
        pixelsStream_s2mPipe_rValid <= pixelsStream_s2mPipe_valid;
      end
      if(pixelsIn_valid) begin
        pixelsIn_rValid <= 1'b1;
      end
      if(pixelsIn_s2mPipe_ready) begin
        pixelsIn_rValid <= 1'b0;
      end
      if(pixelsIn_s2mPipe_ready) begin
        pixelsIn_s2mPipe_rValid <= pixelsIn_s2mPipe_valid;
      end
      if(when_SuperResolutionPart1_l421) begin
        bufferReachRowEnd <= 1'b1;
      end
      if(when_SuperResolutionPart1_l422) begin
        bufferReachFinalRow <= 1'b1;
      end
      if(when_SuperResolutionPart1_l425) begin
        if(bufferReachFinalRow) begin
          bufferReuse <= 1'b1;
          bufferReachRowEnd <= 1'b0;
          bufferReachFinalRow <= 1'b0;
        end else begin
          bufferReachRowEnd <= 1'b0;
        end
      end
      if(when_SuperResolutionPart1_l438) begin
        bufferSwitch <= (! bufferSwitch);
      end
      if(when_SuperResolutionPart1_l439) begin
        holdBuffer <= 1'b1;
        bufferEnable <= 1'b0;
        if(when_SuperResolutionPart1_l442) begin
          writeDone <= 1'b1;
          bufferEnable <= 1'b0;
        end
      end
      if(when_SuperResolutionPart1_l447) begin
        holdBuffer <= 1'b0;
        if(when_SuperResolutionPart1_l449) begin
          nextRowBuffer <= (! nextRowBuffer);
        end
      end
      if(when_SuperResolutionPart1_l453) begin
        frameStart <= 1'b1;
      end
      if(inpDone) begin
        inpDone <= 1'b0;
      end
      controlStateMachine_stateReg <= controlStateMachine_stateNext;
      case(controlStateMachine_stateReg)
        controlStateMachine_enumDef_HOLD : begin
        end
        controlStateMachine_enumDef_PASS : begin
          if(when_SuperResolutionPart1_l507) begin
            frameStart <= 1'b0;
          end
          if(when_SuperResolutionPart1_l510) begin
            outReachRowEnd <= 1'b1;
          end
          if(when_SuperResolutionPart1_l511) begin
            outReachFinalRow <= 1'b1;
          end
          if(when_SuperResolutionPart1_l513) begin
            if(outReachFinalRow) begin
              startRead <= 1'b0;
              readDone <= 1'b1;
              outReachRowEnd <= 1'b0;
              outReachFinalRow <= 1'b0;
            end else begin
              outReachRowEnd <= 1'b0;
            end
          end
          if(controlStream_fire_6) begin
            if(outReachRowEnd) begin
              outReachRowEnd <= 1'b0;
            end
          end
        end
        controlStateMachine_enumDef_ONCE : begin
          if(when_SuperResolutionPart1_l578) begin
            outReachRowEnd <= 1'b1;
          end
          if(when_SuperResolutionPart1_l579) begin
            outReachFinalRow <= 1'b1;
          end
          if(when_SuperResolutionPart1_l581) begin
            if(outReachFinalRow) begin
              startRead <= 1'b0;
              readDone <= 1'b1;
              outReachRowEnd <= 1'b0;
              outReachFinalRow <= 1'b0;
            end else begin
              outReachRowEnd <= 1'b0;
            end
          end
          if(controlStream_fire_12) begin
            if(outReachRowEnd) begin
              outReachRowEnd <= 1'b0;
            end
          end
        end
        controlStateMachine_enumDef_TWICE : begin
          if(when_SuperResolutionPart1_l664) begin
            outReachRowEnd <= 1'b1;
          end
          if(when_SuperResolutionPart1_l665) begin
            outReachFinalRow <= 1'b1;
          end
          if(when_SuperResolutionPart1_l667) begin
            if(outReachFinalRow) begin
              startRead <= 1'b0;
              readDone <= 1'b1;
              outReachRowEnd <= 1'b0;
              outReachFinalRow <= 1'b0;
            end else begin
              outReachRowEnd <= 1'b0;
            end
          end
          if(controlStream_fire_17) begin
            if(outReachRowEnd) begin
              outReachRowEnd <= 1'b0;
            end
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(posedge clk) begin
    startIn_regNext <= startIn;
    if(mainAddrOneStream_ready) begin
      mainAddrOneStream_rData <= mainAddrOneStream_payload;
    end
    if(mainAddrOneStream_s2mPipe_ready) begin
      mainAddrOneStream_s2mPipe_rData <= mainAddrOneStream_s2mPipe_payload;
    end
    if(CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_mainOnePixelStream_payload_1 <= CICC1851_readStage_mainOnePixelStream_payload;
    end
    if(CICC1851_1) begin
      CICC1851_readStage_mainOnePixelStream_payload_2 <= (CICC1851_mainAddrOneStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_mainOnePixelStream_payload_1 : CICC1851_readStage_mainOnePixelStream_payload);
    end
    if(counterAddrOneStream_ready) begin
      counterAddrOneStream_rData <= counterAddrOneStream_payload;
    end
    if(counterAddrOneStream_s2mPipe_ready) begin
      counterAddrOneStream_s2mPipe_rData <= counterAddrOneStream_s2mPipe_payload;
    end
    if(CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_counterOnePixelStream_payload_1 <= CICC1851_readStage_counterOnePixelStream_payload;
    end
    if(CICC1851_2) begin
      CICC1851_readStage_counterOnePixelStream_payload_2 <= (CICC1851_counterAddrOneStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_counterOnePixelStream_payload_1 : CICC1851_readStage_counterOnePixelStream_payload);
    end
    if(mainAddrTwoStream_ready) begin
      mainAddrTwoStream_rData <= mainAddrTwoStream_payload;
    end
    if(mainAddrTwoStream_s2mPipe_ready) begin
      mainAddrTwoStream_s2mPipe_rData <= mainAddrTwoStream_s2mPipe_payload;
    end
    if(CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_mainTwoPixelStream_payload_1 <= CICC1851_readStage_mainTwoPixelStream_payload;
    end
    if(CICC1851_3) begin
      CICC1851_readStage_mainTwoPixelStream_payload_2 <= (CICC1851_mainAddrTwoStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_mainTwoPixelStream_payload_1 : CICC1851_readStage_mainTwoPixelStream_payload);
    end
    if(counterAddrTwoStream_ready) begin
      counterAddrTwoStream_rData <= counterAddrTwoStream_payload;
    end
    if(counterAddrTwoStream_s2mPipe_ready) begin
      counterAddrTwoStream_s2mPipe_rData <= counterAddrTwoStream_s2mPipe_payload;
    end
    if(CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_1) begin
      CICC1851_readStage_counterTwoPixelStream_payload_1 <= CICC1851_readStage_counterTwoPixelStream_payload;
    end
    if(CICC1851_4) begin
      CICC1851_readStage_counterTwoPixelStream_payload_2 <= (CICC1851_counterAddrTwoStream_s2mPipe_m2sPipe_ready_3 ? CICC1851_readStage_counterTwoPixelStream_payload_1 : CICC1851_readStage_counterTwoPixelStream_payload);
    end
    if(controlStream_ready) begin
      controlStream_rData_frameStart <= controlStream_payload_frameStart;
      controlStream_rData_rowEnd <= controlStream_payload_rowEnd;
      controlStream_rData_passMode <= controlStream_payload_passMode;
      controlStream_rData_passValid <= controlStream_payload_passValid;
      controlStream_rData_onceMode <= controlStream_payload_onceMode;
      controlStream_rData_onceValid <= controlStream_payload_onceValid;
      controlStream_rData_mainCompare <= controlStream_payload_mainCompare;
      controlStream_rData_counterCompare <= controlStream_payload_counterCompare;
      controlStream_rData_mainDiff <= controlStream_payload_mainDiff;
      controlStream_rData_counterDiff <= controlStream_payload_counterDiff;
      controlStream_rData_twiceCompValid <= controlStream_payload_twiceCompValid;
      controlStream_rData_twiceMode <= controlStream_payload_twiceMode;
    end
    if(controlStream_s2mPipe_ready) begin
      controlStream_s2mPipe_rData_frameStart <= controlStream_s2mPipe_payload_frameStart;
      controlStream_s2mPipe_rData_rowEnd <= controlStream_s2mPipe_payload_rowEnd;
      controlStream_s2mPipe_rData_passMode <= controlStream_s2mPipe_payload_passMode;
      controlStream_s2mPipe_rData_passValid <= controlStream_s2mPipe_payload_passValid;
      controlStream_s2mPipe_rData_onceMode <= controlStream_s2mPipe_payload_onceMode;
      controlStream_s2mPipe_rData_onceValid <= controlStream_s2mPipe_payload_onceValid;
      controlStream_s2mPipe_rData_mainCompare <= controlStream_s2mPipe_payload_mainCompare;
      controlStream_s2mPipe_rData_counterCompare <= controlStream_s2mPipe_payload_counterCompare;
      controlStream_s2mPipe_rData_mainDiff <= controlStream_s2mPipe_payload_mainDiff;
      controlStream_s2mPipe_rData_counterDiff <= controlStream_s2mPipe_payload_counterDiff;
      controlStream_s2mPipe_rData_twiceCompValid <= controlStream_s2mPipe_payload_twiceCompValid;
      controlStream_s2mPipe_rData_twiceMode <= controlStream_s2mPipe_payload_twiceMode;
    end
    if(controlStream_s2mPipe_m2sPipe_ready) begin
      controlStream_s2mPipe_m2sPipe_rData_frameStart <= controlStream_s2mPipe_m2sPipe_payload_frameStart;
      controlStream_s2mPipe_m2sPipe_rData_rowEnd <= controlStream_s2mPipe_m2sPipe_payload_rowEnd;
      controlStream_s2mPipe_m2sPipe_rData_passMode <= controlStream_s2mPipe_m2sPipe_payload_passMode;
      controlStream_s2mPipe_m2sPipe_rData_passValid <= controlStream_s2mPipe_m2sPipe_payload_passValid;
      controlStream_s2mPipe_m2sPipe_rData_onceMode <= controlStream_s2mPipe_m2sPipe_payload_onceMode;
      controlStream_s2mPipe_m2sPipe_rData_onceValid <= controlStream_s2mPipe_m2sPipe_payload_onceValid;
      controlStream_s2mPipe_m2sPipe_rData_mainCompare <= controlStream_s2mPipe_m2sPipe_payload_mainCompare;
      controlStream_s2mPipe_m2sPipe_rData_counterCompare <= controlStream_s2mPipe_m2sPipe_payload_counterCompare;
      controlStream_s2mPipe_m2sPipe_rData_mainDiff <= controlStream_s2mPipe_m2sPipe_payload_mainDiff;
      controlStream_s2mPipe_m2sPipe_rData_counterDiff <= controlStream_s2mPipe_m2sPipe_payload_counterDiff;
      controlStream_s2mPipe_m2sPipe_rData_twiceCompValid <= controlStream_s2mPipe_m2sPipe_payload_twiceCompValid;
      controlStream_s2mPipe_m2sPipe_rData_twiceMode <= controlStream_s2mPipe_m2sPipe_payload_twiceMode;
    end
    if(controlStream_s2mPipe_m2sPipe_m2sPipe_ready) begin
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_frameStart <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_frameStart;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_rowEnd <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_rowEnd;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_passMode <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passMode;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_passValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_passValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_onceMode <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceMode;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_onceValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_onceValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_mainDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_mainDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_counterDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_counterDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_twiceCompValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceCompValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_rData_twiceMode <= controlStream_s2mPipe_m2sPipe_m2sPipe_payload_twiceMode;
    end
    if(controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_ready) begin
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_frameStart <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_frameStart;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_rowEnd <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_rowEnd;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_passMode <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_passMode;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_passValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_passValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_onceMode <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_onceMode;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_onceValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_onceValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterCompare <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterCompare;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_mainDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_mainDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_counterDiff <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_counterDiff;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_twiceCompValid <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_twiceCompValid;
      controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_rData_twiceMode <= controlStream_s2mPipe_m2sPipe_m2sPipe_s2mPipe_payload_twiceMode;
    end
    if(readStage_mainOnePixelStream_ready) begin
      readStage_mainOnePixelStream_rData <= readStage_mainOnePixelStream_payload;
    end
    if(readStage_mainOnePixelStream_s2mPipe_ready) begin
      readStage_mainOnePixelStream_s2mPipe_rData <= readStage_mainOnePixelStream_s2mPipe_payload;
    end
    if(readStage_counterOnePixelStream_ready) begin
      readStage_counterOnePixelStream_rData <= readStage_counterOnePixelStream_payload;
    end
    if(readStage_counterOnePixelStream_s2mPipe_ready) begin
      readStage_counterOnePixelStream_s2mPipe_rData <= readStage_counterOnePixelStream_s2mPipe_payload;
    end
    if(readStage_mainTwoPixelStream_ready) begin
      readStage_mainTwoPixelStream_rData <= readStage_mainTwoPixelStream_payload;
    end
    if(readStage_mainTwoPixelStream_s2mPipe_ready) begin
      readStage_mainTwoPixelStream_s2mPipe_rData <= readStage_mainTwoPixelStream_s2mPipe_payload;
    end
    if(readStage_counterTwoPixelStream_ready) begin
      readStage_counterTwoPixelStream_rData <= readStage_counterTwoPixelStream_payload;
    end
    if(readStage_counterTwoPixelStream_s2mPipe_ready) begin
      readStage_counterTwoPixelStream_s2mPipe_rData <= readStage_counterTwoPixelStream_s2mPipe_payload;
    end
    if(readStage_controlPipe_translated_ready) begin
      readStage_controlPipe_translated_rData_frameStart <= readStage_controlPipe_translated_payload_frameStart;
      readStage_controlPipe_translated_rData_rowEnd <= readStage_controlPipe_translated_payload_rowEnd;
      readStage_controlPipe_translated_rData_passMode <= readStage_controlPipe_translated_payload_passMode;
      readStage_controlPipe_translated_rData_passValid <= readStage_controlPipe_translated_payload_passValid;
      readStage_controlPipe_translated_rData_onceMode <= readStage_controlPipe_translated_payload_onceMode;
      readStage_controlPipe_translated_rData_onceValid <= readStage_controlPipe_translated_payload_onceValid;
      readStage_controlPipe_translated_rData_mainCompare <= readStage_controlPipe_translated_payload_mainCompare;
      readStage_controlPipe_translated_rData_counterCompare <= readStage_controlPipe_translated_payload_counterCompare;
      readStage_controlPipe_translated_rData_mainDiff <= readStage_controlPipe_translated_payload_mainDiff;
      readStage_controlPipe_translated_rData_counterDiff <= readStage_controlPipe_translated_payload_counterDiff;
      readStage_controlPipe_translated_rData_twiceCompValid <= readStage_controlPipe_translated_payload_twiceCompValid;
      readStage_controlPipe_translated_rData_twiceMode <= readStage_controlPipe_translated_payload_twiceMode;
    end
    if(readStage_controlPipe_translated_s2mPipe_ready) begin
      readStage_controlPipe_translated_s2mPipe_rData_frameStart <= readStage_controlPipe_translated_s2mPipe_payload_frameStart;
      readStage_controlPipe_translated_s2mPipe_rData_rowEnd <= readStage_controlPipe_translated_s2mPipe_payload_rowEnd;
      readStage_controlPipe_translated_s2mPipe_rData_passMode <= readStage_controlPipe_translated_s2mPipe_payload_passMode;
      readStage_controlPipe_translated_s2mPipe_rData_passValid <= readStage_controlPipe_translated_s2mPipe_payload_passValid;
      readStage_controlPipe_translated_s2mPipe_rData_onceMode <= readStage_controlPipe_translated_s2mPipe_payload_onceMode;
      readStage_controlPipe_translated_s2mPipe_rData_onceValid <= readStage_controlPipe_translated_s2mPipe_payload_onceValid;
      readStage_controlPipe_translated_s2mPipe_rData_mainCompare <= readStage_controlPipe_translated_s2mPipe_payload_mainCompare;
      readStage_controlPipe_translated_s2mPipe_rData_counterCompare <= readStage_controlPipe_translated_s2mPipe_payload_counterCompare;
      readStage_controlPipe_translated_s2mPipe_rData_mainDiff <= readStage_controlPipe_translated_s2mPipe_payload_mainDiff;
      readStage_controlPipe_translated_s2mPipe_rData_counterDiff <= readStage_controlPipe_translated_s2mPipe_payload_counterDiff;
      readStage_controlPipe_translated_s2mPipe_rData_twiceCompValid <= readStage_controlPipe_translated_s2mPipe_payload_twiceCompValid;
      readStage_controlPipe_translated_s2mPipe_rData_twiceMode <= readStage_controlPipe_translated_s2mPipe_payload_twiceMode;
    end
    if(compareStage_mainOnePixelStream_ready) begin
      compareStage_mainOnePixelStream_rData <= compareStage_mainOnePixelStream_payload;
    end
    if(compareStage_mainOnePixelStream_s2mPipe_ready) begin
      compareStage_mainOnePixelStream_s2mPipe_rData <= compareStage_mainOnePixelStream_s2mPipe_payload;
    end
    if(compareStage_counterOnePixelStream_ready) begin
      compareStage_counterOnePixelStream_rData <= compareStage_counterOnePixelStream_payload;
    end
    if(compareStage_counterOnePixelStream_s2mPipe_ready) begin
      compareStage_counterOnePixelStream_s2mPipe_rData <= compareStage_counterOnePixelStream_s2mPipe_payload;
    end
    if(compareStage_mainTwoPixelStream_ready) begin
      compareStage_mainTwoPixelStream_rData <= compareStage_mainTwoPixelStream_payload;
    end
    if(compareStage_mainTwoPixelStream_s2mPipe_ready) begin
      compareStage_mainTwoPixelStream_s2mPipe_rData <= compareStage_mainTwoPixelStream_s2mPipe_payload;
    end
    if(compareStage_counterTwoPixelStream_ready) begin
      compareStage_counterTwoPixelStream_rData <= compareStage_counterTwoPixelStream_payload;
    end
    if(compareStage_counterTwoPixelStream_s2mPipe_ready) begin
      compareStage_counterTwoPixelStream_s2mPipe_rData <= compareStage_counterTwoPixelStream_s2mPipe_payload;
    end
    if(compareStage_controlPipe_translated_ready) begin
      compareStage_controlPipe_translated_rData_frameStart <= compareStage_controlPipe_translated_payload_frameStart;
      compareStage_controlPipe_translated_rData_rowEnd <= compareStage_controlPipe_translated_payload_rowEnd;
      compareStage_controlPipe_translated_rData_passMode <= compareStage_controlPipe_translated_payload_passMode;
      compareStage_controlPipe_translated_rData_passValid <= compareStage_controlPipe_translated_payload_passValid;
      compareStage_controlPipe_translated_rData_onceMode <= compareStage_controlPipe_translated_payload_onceMode;
      compareStage_controlPipe_translated_rData_onceValid <= compareStage_controlPipe_translated_payload_onceValid;
      compareStage_controlPipe_translated_rData_mainCompare <= compareStage_controlPipe_translated_payload_mainCompare;
      compareStage_controlPipe_translated_rData_counterCompare <= compareStage_controlPipe_translated_payload_counterCompare;
      compareStage_controlPipe_translated_rData_mainDiff <= compareStage_controlPipe_translated_payload_mainDiff;
      compareStage_controlPipe_translated_rData_counterDiff <= compareStage_controlPipe_translated_payload_counterDiff;
      compareStage_controlPipe_translated_rData_twiceCompValid <= compareStage_controlPipe_translated_payload_twiceCompValid;
      compareStage_controlPipe_translated_rData_twiceMode <= compareStage_controlPipe_translated_payload_twiceMode;
    end
    if(compareStage_controlPipe_translated_s2mPipe_ready) begin
      compareStage_controlPipe_translated_s2mPipe_rData_frameStart <= compareStage_controlPipe_translated_s2mPipe_payload_frameStart;
      compareStage_controlPipe_translated_s2mPipe_rData_rowEnd <= compareStage_controlPipe_translated_s2mPipe_payload_rowEnd;
      compareStage_controlPipe_translated_s2mPipe_rData_passMode <= compareStage_controlPipe_translated_s2mPipe_payload_passMode;
      compareStage_controlPipe_translated_s2mPipe_rData_passValid <= compareStage_controlPipe_translated_s2mPipe_payload_passValid;
      compareStage_controlPipe_translated_s2mPipe_rData_onceMode <= compareStage_controlPipe_translated_s2mPipe_payload_onceMode;
      compareStage_controlPipe_translated_s2mPipe_rData_onceValid <= compareStage_controlPipe_translated_s2mPipe_payload_onceValid;
      compareStage_controlPipe_translated_s2mPipe_rData_mainCompare <= compareStage_controlPipe_translated_s2mPipe_payload_mainCompare;
      compareStage_controlPipe_translated_s2mPipe_rData_counterCompare <= compareStage_controlPipe_translated_s2mPipe_payload_counterCompare;
      compareStage_controlPipe_translated_s2mPipe_rData_mainDiff <= compareStage_controlPipe_translated_s2mPipe_payload_mainDiff;
      compareStage_controlPipe_translated_s2mPipe_rData_counterDiff <= compareStage_controlPipe_translated_s2mPipe_payload_counterDiff;
      compareStage_controlPipe_translated_s2mPipe_rData_twiceCompValid <= compareStage_controlPipe_translated_s2mPipe_payload_twiceCompValid;
      compareStage_controlPipe_translated_s2mPipe_rData_twiceMode <= compareStage_controlPipe_translated_s2mPipe_payload_twiceMode;
    end
    if(diffStage_mainOnePixelStream_ready) begin
      diffStage_mainOnePixelStream_rData <= diffStage_mainOnePixelStream_payload;
    end
    if(diffStage_mainOnePixelStream_s2mPipe_ready) begin
      diffStage_mainOnePixelStream_s2mPipe_rData <= diffStage_mainOnePixelStream_s2mPipe_payload;
    end
    if(diffStage_counterOnePixelStream_ready) begin
      diffStage_counterOnePixelStream_rData <= diffStage_counterOnePixelStream_payload;
    end
    if(diffStage_counterOnePixelStream_s2mPipe_ready) begin
      diffStage_counterOnePixelStream_s2mPipe_rData <= diffStage_counterOnePixelStream_s2mPipe_payload;
    end
    if(diffStage_mainTwoPixelStream_ready) begin
      diffStage_mainTwoPixelStream_rData <= diffStage_mainTwoPixelStream_payload;
    end
    if(diffStage_mainTwoPixelStream_s2mPipe_ready) begin
      diffStage_mainTwoPixelStream_s2mPipe_rData <= diffStage_mainTwoPixelStream_s2mPipe_payload;
    end
    if(diffStage_counterTwoPixelStream_ready) begin
      diffStage_counterTwoPixelStream_rData <= diffStage_counterTwoPixelStream_payload;
    end
    if(diffStage_counterTwoPixelStream_s2mPipe_ready) begin
      diffStage_counterTwoPixelStream_s2mPipe_rData <= diffStage_counterTwoPixelStream_s2mPipe_payload;
    end
    if(diffStage_controlPipe_fork_io_outputs_0_ready) begin
      diffStage_controlPipe_fork_io_outputs_0_rData_frameStart <= diffStage_controlPipe_fork_io_outputs_0_payload_frameStart;
      diffStage_controlPipe_fork_io_outputs_0_rData_rowEnd <= diffStage_controlPipe_fork_io_outputs_0_payload_rowEnd;
      diffStage_controlPipe_fork_io_outputs_0_rData_passMode <= diffStage_controlPipe_fork_io_outputs_0_payload_passMode;
      diffStage_controlPipe_fork_io_outputs_0_rData_passValid <= diffStage_controlPipe_fork_io_outputs_0_payload_passValid;
      diffStage_controlPipe_fork_io_outputs_0_rData_onceMode <= diffStage_controlPipe_fork_io_outputs_0_payload_onceMode;
      diffStage_controlPipe_fork_io_outputs_0_rData_onceValid <= diffStage_controlPipe_fork_io_outputs_0_payload_onceValid;
      diffStage_controlPipe_fork_io_outputs_0_rData_mainCompare <= diffStage_controlPipe_fork_io_outputs_0_payload_mainCompare;
      diffStage_controlPipe_fork_io_outputs_0_rData_counterCompare <= diffStage_controlPipe_fork_io_outputs_0_payload_counterCompare;
      diffStage_controlPipe_fork_io_outputs_0_rData_mainDiff <= diffStage_controlPipe_fork_io_outputs_0_payload_mainDiff;
      diffStage_controlPipe_fork_io_outputs_0_rData_counterDiff <= diffStage_controlPipe_fork_io_outputs_0_payload_counterDiff;
      diffStage_controlPipe_fork_io_outputs_0_rData_twiceCompValid <= diffStage_controlPipe_fork_io_outputs_0_payload_twiceCompValid;
      diffStage_controlPipe_fork_io_outputs_0_rData_twiceMode <= diffStage_controlPipe_fork_io_outputs_0_payload_twiceMode;
    end
    if(diffStage_controlPipe_fork_io_outputs_0_s2mPipe_ready) begin
      diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_frameStart <= diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_frameStart;
      diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_rowEnd <= diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_rowEnd;
      diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_passMode <= diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_passMode;
      diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_passValid <= diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_passValid;
      diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_onceMode <= diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_onceMode;
      diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_onceValid <= diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_onceValid;
      diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_mainCompare <= diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_mainCompare;
      diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_counterCompare <= diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_counterCompare;
      diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_mainDiff <= diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_mainDiff;
      diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_counterDiff <= diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_counterDiff;
      diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_twiceCompValid <= diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_twiceCompValid;
      diffStage_controlPipe_fork_io_outputs_0_s2mPipe_rData_twiceMode <= diffStage_controlPipe_fork_io_outputs_0_s2mPipe_payload_twiceMode;
    end
    if(resultStage_pixelStream_ready) begin
      resultStage_pixelStream_rData <= resultStage_pixelStream_payload;
    end
    if(resultStage_pixelStream_s2mPipe_ready) begin
      resultStage_pixelStream_s2mPipe_rData <= resultStage_pixelStream_s2mPipe_payload;
    end
    if(pixelsStream_ready) begin
      pixelsStream_rData_pixel <= pixelsStream_payload_pixel;
      pixelsStream_rData_frameStart <= pixelsStream_payload_frameStart;
      pixelsStream_rData_rowEnd <= pixelsStream_payload_rowEnd;
    end
    if(pixelsStream_s2mPipe_ready) begin
      pixelsStream_s2mPipe_rData_pixel <= pixelsStream_s2mPipe_payload_pixel;
      pixelsStream_s2mPipe_rData_frameStart <= pixelsStream_s2mPipe_payload_frameStart;
      pixelsStream_s2mPipe_rData_rowEnd <= pixelsStream_s2mPipe_payload_rowEnd;
    end
    if(pixelsIn_ready) begin
      pixelsIn_rData_pixel <= pixelsIn_payload_pixel;
      pixelsIn_rData_frameStart <= pixelsIn_payload_frameStart;
      pixelsIn_rData_rowEnd <= pixelsIn_payload_rowEnd;
    end
    if(pixelsIn_s2mPipe_ready) begin
      pixelsIn_s2mPipe_rData_pixel <= pixelsIn_s2mPipe_payload_pixel;
      pixelsIn_s2mPipe_rData_frameStart <= pixelsIn_s2mPipe_payload_frameStart;
      pixelsIn_s2mPipe_rData_rowEnd <= pixelsIn_s2mPipe_payload_rowEnd;
    end
  end


endmodule

module ChannelMasterTransformer (
  input               allPixelChannelIn_valid,
  output              allPixelChannelIn_ready,
  input      [31:0]   allPixelChannelIn_payload_pixel,
  input               allPixelChannelIn_payload_frameStart,
  input               allPixelChannelIn_payload_rowEnd,
  output              bPixelChannelOut_valid,
  input               bPixelChannelOut_ready,
  output     [7:0]    bPixelChannelOut_payload_pixel,
  output              bPixelChannelOut_payload_frameStart,
  output              bPixelChannelOut_payload_rowEnd,
  output              gPixelChannelOut_valid,
  input               gPixelChannelOut_ready,
  output     [7:0]    gPixelChannelOut_payload_pixel,
  output              gPixelChannelOut_payload_frameStart,
  output              gPixelChannelOut_payload_rowEnd,
  output              rPixelChannelOut_valid,
  input               rPixelChannelOut_ready,
  output     [7:0]    rPixelChannelOut_payload_pixel,
  output              rPixelChannelOut_payload_frameStart,
  output              rPixelChannelOut_payload_rowEnd,
  input               clk,
  input               resetn
);

  wire                allPixelChannelIn_fork_io_input_ready;
  wire                allPixelChannelIn_fork_io_outputs_0_valid;
  wire       [31:0]   allPixelChannelIn_fork_io_outputs_0_payload_pixel;
  wire                allPixelChannelIn_fork_io_outputs_0_payload_frameStart;
  wire                allPixelChannelIn_fork_io_outputs_0_payload_rowEnd;
  wire                allPixelChannelIn_fork_io_outputs_1_valid;
  wire       [31:0]   allPixelChannelIn_fork_io_outputs_1_payload_pixel;
  wire                allPixelChannelIn_fork_io_outputs_1_payload_frameStart;
  wire                allPixelChannelIn_fork_io_outputs_1_payload_rowEnd;
  wire                allPixelChannelIn_fork_io_outputs_2_valid;
  wire       [31:0]   allPixelChannelIn_fork_io_outputs_2_payload_pixel;
  wire                allPixelChannelIn_fork_io_outputs_2_payload_frameStart;
  wire                allPixelChannelIn_fork_io_outputs_2_payload_rowEnd;
  wire                allPixelChannelIn_fork_io_outputs_0_translated_valid;
  wire                allPixelChannelIn_fork_io_outputs_0_translated_ready;
  wire       [7:0]    allPixelChannelIn_fork_io_outputs_0_translated_payload_pixel;
  wire                allPixelChannelIn_fork_io_outputs_0_translated_payload_frameStart;
  wire                allPixelChannelIn_fork_io_outputs_0_translated_payload_rowEnd;
  wire                allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_valid;
  reg                 allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_ready;
  wire       [7:0]    allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_payload_pixel;
  wire                allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_payload_frameStart;
  wire                allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_payload_rowEnd;
  reg                 allPixelChannelIn_fork_io_outputs_0_translated_rValid;
  reg        [7:0]    allPixelChannelIn_fork_io_outputs_0_translated_rData_pixel;
  reg                 allPixelChannelIn_fork_io_outputs_0_translated_rData_frameStart;
  reg                 allPixelChannelIn_fork_io_outputs_0_translated_rData_rowEnd;
  wire                allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_m2sPipe_valid;
  wire                allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_m2sPipe_ready;
  wire       [7:0]    allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_m2sPipe_payload_pixel;
  wire                allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_m2sPipe_payload_frameStart;
  wire                allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_m2sPipe_payload_rowEnd;
  reg                 allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_rValid;
  reg        [7:0]    allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_rData_pixel;
  reg                 allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_rData_frameStart;
  reg                 allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_rData_rowEnd;
  wire                when_Stream_l368;
  wire                allPixelChannelIn_fork_io_outputs_1_translated_valid;
  wire                allPixelChannelIn_fork_io_outputs_1_translated_ready;
  wire       [7:0]    allPixelChannelIn_fork_io_outputs_1_translated_payload_pixel;
  wire                allPixelChannelIn_fork_io_outputs_1_translated_payload_frameStart;
  wire                allPixelChannelIn_fork_io_outputs_1_translated_payload_rowEnd;
  wire                allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_valid;
  reg                 allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_ready;
  wire       [7:0]    allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_payload_pixel;
  wire                allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_payload_frameStart;
  wire                allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_payload_rowEnd;
  reg                 allPixelChannelIn_fork_io_outputs_1_translated_rValid;
  reg        [7:0]    allPixelChannelIn_fork_io_outputs_1_translated_rData_pixel;
  reg                 allPixelChannelIn_fork_io_outputs_1_translated_rData_frameStart;
  reg                 allPixelChannelIn_fork_io_outputs_1_translated_rData_rowEnd;
  wire                allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_m2sPipe_valid;
  wire                allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_m2sPipe_ready;
  wire       [7:0]    allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_m2sPipe_payload_pixel;
  wire                allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_m2sPipe_payload_frameStart;
  wire                allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_m2sPipe_payload_rowEnd;
  reg                 allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_rValid;
  reg        [7:0]    allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_rData_pixel;
  reg                 allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_rData_frameStart;
  reg                 allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_rData_rowEnd;
  wire                when_Stream_l368_1;
  wire                allPixelChannelIn_fork_io_outputs_2_translated_valid;
  wire                allPixelChannelIn_fork_io_outputs_2_translated_ready;
  wire       [7:0]    allPixelChannelIn_fork_io_outputs_2_translated_payload_pixel;
  wire                allPixelChannelIn_fork_io_outputs_2_translated_payload_frameStart;
  wire                allPixelChannelIn_fork_io_outputs_2_translated_payload_rowEnd;
  wire                allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_valid;
  reg                 allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_ready;
  wire       [7:0]    allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_payload_pixel;
  wire                allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_payload_frameStart;
  wire                allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_payload_rowEnd;
  reg                 allPixelChannelIn_fork_io_outputs_2_translated_rValid;
  reg        [7:0]    allPixelChannelIn_fork_io_outputs_2_translated_rData_pixel;
  reg                 allPixelChannelIn_fork_io_outputs_2_translated_rData_frameStart;
  reg                 allPixelChannelIn_fork_io_outputs_2_translated_rData_rowEnd;
  wire                allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_m2sPipe_valid;
  wire                allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_m2sPipe_ready;
  wire       [7:0]    allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_m2sPipe_payload_pixel;
  wire                allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_m2sPipe_payload_frameStart;
  wire                allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_m2sPipe_payload_rowEnd;
  reg                 allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_rValid;
  reg        [7:0]    allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_rData_pixel;
  reg                 allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_rData_frameStart;
  reg                 allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_rData_rowEnd;
  wire                when_Stream_l368_2;

  StreamFork allPixelChannelIn_fork (
    .io_input_valid                  (allPixelChannelIn_valid                                ), //i
    .io_input_ready                  (allPixelChannelIn_fork_io_input_ready                  ), //o
    .io_input_payload_pixel          (allPixelChannelIn_payload_pixel[31:0]                  ), //i
    .io_input_payload_frameStart     (allPixelChannelIn_payload_frameStart                   ), //i
    .io_input_payload_rowEnd         (allPixelChannelIn_payload_rowEnd                       ), //i
    .io_outputs_0_valid              (allPixelChannelIn_fork_io_outputs_0_valid              ), //o
    .io_outputs_0_ready              (allPixelChannelIn_fork_io_outputs_0_translated_ready   ), //i
    .io_outputs_0_payload_pixel      (allPixelChannelIn_fork_io_outputs_0_payload_pixel[31:0]), //o
    .io_outputs_0_payload_frameStart (allPixelChannelIn_fork_io_outputs_0_payload_frameStart ), //o
    .io_outputs_0_payload_rowEnd     (allPixelChannelIn_fork_io_outputs_0_payload_rowEnd     ), //o
    .io_outputs_1_valid              (allPixelChannelIn_fork_io_outputs_1_valid              ), //o
    .io_outputs_1_ready              (allPixelChannelIn_fork_io_outputs_1_translated_ready   ), //i
    .io_outputs_1_payload_pixel      (allPixelChannelIn_fork_io_outputs_1_payload_pixel[31:0]), //o
    .io_outputs_1_payload_frameStart (allPixelChannelIn_fork_io_outputs_1_payload_frameStart ), //o
    .io_outputs_1_payload_rowEnd     (allPixelChannelIn_fork_io_outputs_1_payload_rowEnd     ), //o
    .io_outputs_2_valid              (allPixelChannelIn_fork_io_outputs_2_valid              ), //o
    .io_outputs_2_ready              (allPixelChannelIn_fork_io_outputs_2_translated_ready   ), //i
    .io_outputs_2_payload_pixel      (allPixelChannelIn_fork_io_outputs_2_payload_pixel[31:0]), //o
    .io_outputs_2_payload_frameStart (allPixelChannelIn_fork_io_outputs_2_payload_frameStart ), //o
    .io_outputs_2_payload_rowEnd     (allPixelChannelIn_fork_io_outputs_2_payload_rowEnd     )  //o
  );
  assign allPixelChannelIn_ready = allPixelChannelIn_fork_io_input_ready;
  assign allPixelChannelIn_fork_io_outputs_0_translated_valid = allPixelChannelIn_fork_io_outputs_0_valid;
  assign allPixelChannelIn_fork_io_outputs_0_translated_payload_pixel = allPixelChannelIn_fork_io_outputs_0_payload_pixel[7 : 0];
  assign allPixelChannelIn_fork_io_outputs_0_translated_payload_frameStart = allPixelChannelIn_fork_io_outputs_0_payload_frameStart;
  assign allPixelChannelIn_fork_io_outputs_0_translated_payload_rowEnd = allPixelChannelIn_fork_io_outputs_0_payload_rowEnd;
  assign allPixelChannelIn_fork_io_outputs_0_translated_ready = (! allPixelChannelIn_fork_io_outputs_0_translated_rValid);
  assign allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_valid = (allPixelChannelIn_fork_io_outputs_0_translated_valid || allPixelChannelIn_fork_io_outputs_0_translated_rValid);
  assign allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_payload_pixel = (allPixelChannelIn_fork_io_outputs_0_translated_rValid ? allPixelChannelIn_fork_io_outputs_0_translated_rData_pixel : allPixelChannelIn_fork_io_outputs_0_translated_payload_pixel);
  assign allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_payload_frameStart = (allPixelChannelIn_fork_io_outputs_0_translated_rValid ? allPixelChannelIn_fork_io_outputs_0_translated_rData_frameStart : allPixelChannelIn_fork_io_outputs_0_translated_payload_frameStart);
  assign allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_payload_rowEnd = (allPixelChannelIn_fork_io_outputs_0_translated_rValid ? allPixelChannelIn_fork_io_outputs_0_translated_rData_rowEnd : allPixelChannelIn_fork_io_outputs_0_translated_payload_rowEnd);
  always @(*) begin
    allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_ready = allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368) begin
      allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368 = (! allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_m2sPipe_valid);
  assign allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_m2sPipe_valid = allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_rValid;
  assign allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_m2sPipe_payload_pixel = allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_rData_pixel;
  assign allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_m2sPipe_payload_frameStart = allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_rData_frameStart;
  assign allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_m2sPipe_payload_rowEnd = allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_rData_rowEnd;
  assign bPixelChannelOut_valid = allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_m2sPipe_valid;
  assign allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_m2sPipe_ready = bPixelChannelOut_ready;
  assign bPixelChannelOut_payload_pixel = allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_m2sPipe_payload_pixel;
  assign bPixelChannelOut_payload_frameStart = allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_m2sPipe_payload_frameStart;
  assign bPixelChannelOut_payload_rowEnd = allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_m2sPipe_payload_rowEnd;
  assign allPixelChannelIn_fork_io_outputs_1_translated_valid = allPixelChannelIn_fork_io_outputs_1_valid;
  assign allPixelChannelIn_fork_io_outputs_1_translated_payload_pixel = allPixelChannelIn_fork_io_outputs_1_payload_pixel[15 : 8];
  assign allPixelChannelIn_fork_io_outputs_1_translated_payload_frameStart = allPixelChannelIn_fork_io_outputs_1_payload_frameStart;
  assign allPixelChannelIn_fork_io_outputs_1_translated_payload_rowEnd = allPixelChannelIn_fork_io_outputs_1_payload_rowEnd;
  assign allPixelChannelIn_fork_io_outputs_1_translated_ready = (! allPixelChannelIn_fork_io_outputs_1_translated_rValid);
  assign allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_valid = (allPixelChannelIn_fork_io_outputs_1_translated_valid || allPixelChannelIn_fork_io_outputs_1_translated_rValid);
  assign allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_payload_pixel = (allPixelChannelIn_fork_io_outputs_1_translated_rValid ? allPixelChannelIn_fork_io_outputs_1_translated_rData_pixel : allPixelChannelIn_fork_io_outputs_1_translated_payload_pixel);
  assign allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_payload_frameStart = (allPixelChannelIn_fork_io_outputs_1_translated_rValid ? allPixelChannelIn_fork_io_outputs_1_translated_rData_frameStart : allPixelChannelIn_fork_io_outputs_1_translated_payload_frameStart);
  assign allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_payload_rowEnd = (allPixelChannelIn_fork_io_outputs_1_translated_rValid ? allPixelChannelIn_fork_io_outputs_1_translated_rData_rowEnd : allPixelChannelIn_fork_io_outputs_1_translated_payload_rowEnd);
  always @(*) begin
    allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_ready = allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_1) begin
      allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_1 = (! allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_m2sPipe_valid);
  assign allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_m2sPipe_valid = allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_rValid;
  assign allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_m2sPipe_payload_pixel = allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_rData_pixel;
  assign allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_m2sPipe_payload_frameStart = allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_rData_frameStart;
  assign allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_m2sPipe_payload_rowEnd = allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_rData_rowEnd;
  assign gPixelChannelOut_valid = allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_m2sPipe_valid;
  assign allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_m2sPipe_ready = gPixelChannelOut_ready;
  assign gPixelChannelOut_payload_pixel = allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_m2sPipe_payload_pixel;
  assign gPixelChannelOut_payload_frameStart = allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_m2sPipe_payload_frameStart;
  assign gPixelChannelOut_payload_rowEnd = allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_m2sPipe_payload_rowEnd;
  assign allPixelChannelIn_fork_io_outputs_2_translated_valid = allPixelChannelIn_fork_io_outputs_2_valid;
  assign allPixelChannelIn_fork_io_outputs_2_translated_payload_pixel = allPixelChannelIn_fork_io_outputs_2_payload_pixel[23 : 16];
  assign allPixelChannelIn_fork_io_outputs_2_translated_payload_frameStart = allPixelChannelIn_fork_io_outputs_2_payload_frameStart;
  assign allPixelChannelIn_fork_io_outputs_2_translated_payload_rowEnd = allPixelChannelIn_fork_io_outputs_2_payload_rowEnd;
  assign allPixelChannelIn_fork_io_outputs_2_translated_ready = (! allPixelChannelIn_fork_io_outputs_2_translated_rValid);
  assign allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_valid = (allPixelChannelIn_fork_io_outputs_2_translated_valid || allPixelChannelIn_fork_io_outputs_2_translated_rValid);
  assign allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_payload_pixel = (allPixelChannelIn_fork_io_outputs_2_translated_rValid ? allPixelChannelIn_fork_io_outputs_2_translated_rData_pixel : allPixelChannelIn_fork_io_outputs_2_translated_payload_pixel);
  assign allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_payload_frameStart = (allPixelChannelIn_fork_io_outputs_2_translated_rValid ? allPixelChannelIn_fork_io_outputs_2_translated_rData_frameStart : allPixelChannelIn_fork_io_outputs_2_translated_payload_frameStart);
  assign allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_payload_rowEnd = (allPixelChannelIn_fork_io_outputs_2_translated_rValid ? allPixelChannelIn_fork_io_outputs_2_translated_rData_rowEnd : allPixelChannelIn_fork_io_outputs_2_translated_payload_rowEnd);
  always @(*) begin
    allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_ready = allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_2) begin
      allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_2 = (! allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_m2sPipe_valid);
  assign allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_m2sPipe_valid = allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_rValid;
  assign allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_m2sPipe_payload_pixel = allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_rData_pixel;
  assign allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_m2sPipe_payload_frameStart = allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_rData_frameStart;
  assign allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_m2sPipe_payload_rowEnd = allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_rData_rowEnd;
  assign rPixelChannelOut_valid = allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_m2sPipe_valid;
  assign allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_m2sPipe_ready = rPixelChannelOut_ready;
  assign rPixelChannelOut_payload_pixel = allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_m2sPipe_payload_pixel;
  assign rPixelChannelOut_payload_frameStart = allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_m2sPipe_payload_frameStart;
  assign rPixelChannelOut_payload_rowEnd = allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_m2sPipe_payload_rowEnd;
  always @(posedge clk or negedge resetn) begin
    if(!resetn) begin
      allPixelChannelIn_fork_io_outputs_0_translated_rValid <= 1'b0;
      allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_rValid <= 1'b0;
      allPixelChannelIn_fork_io_outputs_1_translated_rValid <= 1'b0;
      allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_rValid <= 1'b0;
      allPixelChannelIn_fork_io_outputs_2_translated_rValid <= 1'b0;
      allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_rValid <= 1'b0;
    end else begin
      if(allPixelChannelIn_fork_io_outputs_0_translated_valid) begin
        allPixelChannelIn_fork_io_outputs_0_translated_rValid <= 1'b1;
      end
      if(allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_ready) begin
        allPixelChannelIn_fork_io_outputs_0_translated_rValid <= 1'b0;
      end
      if(allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_ready) begin
        allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_rValid <= allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_valid;
      end
      if(allPixelChannelIn_fork_io_outputs_1_translated_valid) begin
        allPixelChannelIn_fork_io_outputs_1_translated_rValid <= 1'b1;
      end
      if(allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_ready) begin
        allPixelChannelIn_fork_io_outputs_1_translated_rValid <= 1'b0;
      end
      if(allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_ready) begin
        allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_rValid <= allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_valid;
      end
      if(allPixelChannelIn_fork_io_outputs_2_translated_valid) begin
        allPixelChannelIn_fork_io_outputs_2_translated_rValid <= 1'b1;
      end
      if(allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_ready) begin
        allPixelChannelIn_fork_io_outputs_2_translated_rValid <= 1'b0;
      end
      if(allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_ready) begin
        allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_rValid <= allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_valid;
      end
    end
  end

  always @(posedge clk) begin
    if(allPixelChannelIn_fork_io_outputs_0_translated_ready) begin
      allPixelChannelIn_fork_io_outputs_0_translated_rData_pixel <= allPixelChannelIn_fork_io_outputs_0_translated_payload_pixel;
      allPixelChannelIn_fork_io_outputs_0_translated_rData_frameStart <= allPixelChannelIn_fork_io_outputs_0_translated_payload_frameStart;
      allPixelChannelIn_fork_io_outputs_0_translated_rData_rowEnd <= allPixelChannelIn_fork_io_outputs_0_translated_payload_rowEnd;
    end
    if(allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_ready) begin
      allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_rData_pixel <= allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_payload_pixel;
      allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_rData_frameStart <= allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_payload_frameStart;
      allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_rData_rowEnd <= allPixelChannelIn_fork_io_outputs_0_translated_s2mPipe_payload_rowEnd;
    end
    if(allPixelChannelIn_fork_io_outputs_1_translated_ready) begin
      allPixelChannelIn_fork_io_outputs_1_translated_rData_pixel <= allPixelChannelIn_fork_io_outputs_1_translated_payload_pixel;
      allPixelChannelIn_fork_io_outputs_1_translated_rData_frameStart <= allPixelChannelIn_fork_io_outputs_1_translated_payload_frameStart;
      allPixelChannelIn_fork_io_outputs_1_translated_rData_rowEnd <= allPixelChannelIn_fork_io_outputs_1_translated_payload_rowEnd;
    end
    if(allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_ready) begin
      allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_rData_pixel <= allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_payload_pixel;
      allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_rData_frameStart <= allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_payload_frameStart;
      allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_rData_rowEnd <= allPixelChannelIn_fork_io_outputs_1_translated_s2mPipe_payload_rowEnd;
    end
    if(allPixelChannelIn_fork_io_outputs_2_translated_ready) begin
      allPixelChannelIn_fork_io_outputs_2_translated_rData_pixel <= allPixelChannelIn_fork_io_outputs_2_translated_payload_pixel;
      allPixelChannelIn_fork_io_outputs_2_translated_rData_frameStart <= allPixelChannelIn_fork_io_outputs_2_translated_payload_frameStart;
      allPixelChannelIn_fork_io_outputs_2_translated_rData_rowEnd <= allPixelChannelIn_fork_io_outputs_2_translated_payload_rowEnd;
    end
    if(allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_ready) begin
      allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_rData_pixel <= allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_payload_pixel;
      allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_rData_frameStart <= allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_payload_frameStart;
      allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_rData_rowEnd <= allPixelChannelIn_fork_io_outputs_2_translated_s2mPipe_payload_rowEnd;
    end
  end


endmodule

module DDRDataWrapper (
  input               ddrIn_valid,
  output reg          ddrIn_ready,
  input      [31:0]   ddrIn_payload,
  output              pixelsOut_valid,
  input               pixelsOut_ready,
  output     [31:0]   pixelsOut_payload_pixel,
  output              pixelsOut_payload_frameStart,
  output              pixelsOut_payload_rowEnd,
  input               inpDone,
  input      [9:0]    bmpWidth,
  input               clk,
  input               resetn
);

  wire       [9:0]    transactionCounter_io_count;
  wire                transactionCounter_io_working;
  wire                transactionCounter_io_last;
  wire                transactionCounter_io_done;
  wire       [9:0]    transactionCounter_io_value;
  reg                 isNewTransfer;
  wire                pixelsOut_fire;
  wire                when_DDRDataWrapper_l20;
  reg        [9:0]    imgWidth;
  wire                ddrIn_fire;
  wire                pixelsOut_fire_1;
  wire                ddrIn_m2sPipe_valid;
  wire                ddrIn_m2sPipe_ready;
  wire       [31:0]   ddrIn_m2sPipe_payload;
  reg                 ddrIn_rValid;
  reg        [31:0]   ddrIn_rData;
  wire                when_Stream_l368;

  StreamTransactionCounter transactionCounter (
    .io_ctrlFire   (ddrIn_fire                      ), //i
    .io_targetFire (pixelsOut_fire_1                ), //i
    .io_count      (transactionCounter_io_count[9:0]), //i
    .io_working    (transactionCounter_io_working   ), //o
    .io_last       (transactionCounter_io_last      ), //o
    .io_done       (transactionCounter_io_done      ), //o
    .io_value      (transactionCounter_io_value[9:0]), //o
    .clk           (clk                             ), //i
    .resetn        (resetn                          )  //i
  );
  assign pixelsOut_fire = (pixelsOut_valid && pixelsOut_ready);
  assign when_DDRDataWrapper_l20 = (pixelsOut_payload_frameStart && pixelsOut_fire);
  assign ddrIn_fire = (ddrIn_valid && ddrIn_ready);
  assign pixelsOut_fire_1 = (pixelsOut_valid && pixelsOut_ready);
  assign transactionCounter_io_count = (imgWidth - 10'h001);
  always @(*) begin
    ddrIn_ready = ddrIn_m2sPipe_ready;
    if(when_Stream_l368) begin
      ddrIn_ready = 1'b1;
    end
  end

  assign when_Stream_l368 = (! ddrIn_m2sPipe_valid);
  assign ddrIn_m2sPipe_valid = ddrIn_rValid;
  assign ddrIn_m2sPipe_payload = ddrIn_rData;
  assign pixelsOut_valid = ddrIn_m2sPipe_valid;
  assign ddrIn_m2sPipe_ready = pixelsOut_ready;
  assign pixelsOut_payload_pixel = ddrIn_m2sPipe_payload;
  assign pixelsOut_payload_rowEnd = transactionCounter_io_last;
  assign pixelsOut_payload_frameStart = (isNewTransfer && (transactionCounter_io_value == 10'h0));
  always @(posedge clk or negedge resetn) begin
    if(!resetn) begin
      isNewTransfer <= 1'b1;
      imgWidth <= 10'h3ff;
      ddrIn_rValid <= 1'b0;
    end else begin
      if(inpDone) begin
        isNewTransfer <= 1'b1;
      end
      if(when_DDRDataWrapper_l20) begin
        isNewTransfer <= 1'b0;
      end
      imgWidth <= bmpWidth;
      if(ddrIn_ready) begin
        ddrIn_rValid <= ddrIn_valid;
      end
    end
  end

  always @(posedge clk) begin
    if(ddrIn_ready) begin
      ddrIn_rData <= ddrIn_payload;
    end
  end


endmodule

//StreamFork_3 replaced by StreamFork_3

//StreamFork_2 replaced by StreamFork_2

//StreamFork_1 replaced by StreamFork_1

//StreamFork_3 replaced by StreamFork_3

//StreamFork_2 replaced by StreamFork_2

//StreamFork_1 replaced by StreamFork_1

module StreamFork_3 (
  input               io_input_valid,
  output              io_input_ready,
  input               io_input_payload_frameStart,
  input               io_input_payload_rowEnd,
  input               io_input_payload_pipeValid,
  input               io_input_payload_firstRow,
  input               io_input_payload_lastRow,
  input               io_input_payload_finalResult,
  input               io_input_payload_mainCompare,
  input               io_input_payload_counterCompare,
  input               io_input_payload_horizontalCompare,
  input               io_input_payload_verticalCompare,
  input      [7:0]    io_input_payload_mainDiff,
  input      [7:0]    io_input_payload_counterDiff,
  input      [7:0]    io_input_payload_horizontalDiff,
  input      [7:0]    io_input_payload_verticalDiff,
  input               io_input_payload_isHorizontalMin,
  input      [7:0]    io_input_payload_minDiff,
  input      [1:0]    io_input_payload_currentPosition,
  input      [1:0]    io_input_payload_nextPosition,
  input               io_input_payload_horizontalDirectionValid,
  input               io_input_payload_verticalDirectionValid,
  input               io_input_payload_mainDirectionValid,
  input               io_input_payload_counterDirectionValid,
  input               io_input_payload_inValidMinDiff,
  output              io_outputs_0_valid,
  input               io_outputs_0_ready,
  output              io_outputs_0_payload_frameStart,
  output              io_outputs_0_payload_rowEnd,
  output              io_outputs_0_payload_pipeValid,
  output              io_outputs_0_payload_firstRow,
  output              io_outputs_0_payload_lastRow,
  output              io_outputs_0_payload_finalResult,
  output              io_outputs_0_payload_mainCompare,
  output              io_outputs_0_payload_counterCompare,
  output              io_outputs_0_payload_horizontalCompare,
  output              io_outputs_0_payload_verticalCompare,
  output     [7:0]    io_outputs_0_payload_mainDiff,
  output     [7:0]    io_outputs_0_payload_counterDiff,
  output     [7:0]    io_outputs_0_payload_horizontalDiff,
  output     [7:0]    io_outputs_0_payload_verticalDiff,
  output              io_outputs_0_payload_isHorizontalMin,
  output     [7:0]    io_outputs_0_payload_minDiff,
  output     [1:0]    io_outputs_0_payload_currentPosition,
  output     [1:0]    io_outputs_0_payload_nextPosition,
  output              io_outputs_0_payload_horizontalDirectionValid,
  output              io_outputs_0_payload_verticalDirectionValid,
  output              io_outputs_0_payload_mainDirectionValid,
  output              io_outputs_0_payload_counterDirectionValid,
  output              io_outputs_0_payload_inValidMinDiff,
  output              io_outputs_1_valid,
  input               io_outputs_1_ready,
  output              io_outputs_1_payload_frameStart,
  output              io_outputs_1_payload_rowEnd,
  output              io_outputs_1_payload_pipeValid,
  output              io_outputs_1_payload_firstRow,
  output              io_outputs_1_payload_lastRow,
  output              io_outputs_1_payload_finalResult,
  output              io_outputs_1_payload_mainCompare,
  output              io_outputs_1_payload_counterCompare,
  output              io_outputs_1_payload_horizontalCompare,
  output              io_outputs_1_payload_verticalCompare,
  output     [7:0]    io_outputs_1_payload_mainDiff,
  output     [7:0]    io_outputs_1_payload_counterDiff,
  output     [7:0]    io_outputs_1_payload_horizontalDiff,
  output     [7:0]    io_outputs_1_payload_verticalDiff,
  output              io_outputs_1_payload_isHorizontalMin,
  output     [7:0]    io_outputs_1_payload_minDiff,
  output     [1:0]    io_outputs_1_payload_currentPosition,
  output     [1:0]    io_outputs_1_payload_nextPosition,
  output              io_outputs_1_payload_horizontalDirectionValid,
  output              io_outputs_1_payload_verticalDirectionValid,
  output              io_outputs_1_payload_mainDirectionValid,
  output              io_outputs_1_payload_counterDirectionValid,
  output              io_outputs_1_payload_inValidMinDiff
);


  assign io_input_ready = (io_outputs_0_ready && io_outputs_1_ready);
  assign io_outputs_0_valid = (io_input_valid && io_input_ready);
  assign io_outputs_1_valid = (io_input_valid && io_input_ready);
  assign io_outputs_0_payload_frameStart = io_input_payload_frameStart;
  assign io_outputs_0_payload_rowEnd = io_input_payload_rowEnd;
  assign io_outputs_0_payload_pipeValid = io_input_payload_pipeValid;
  assign io_outputs_0_payload_firstRow = io_input_payload_firstRow;
  assign io_outputs_0_payload_lastRow = io_input_payload_lastRow;
  assign io_outputs_0_payload_finalResult = io_input_payload_finalResult;
  assign io_outputs_0_payload_mainCompare = io_input_payload_mainCompare;
  assign io_outputs_0_payload_counterCompare = io_input_payload_counterCompare;
  assign io_outputs_0_payload_horizontalCompare = io_input_payload_horizontalCompare;
  assign io_outputs_0_payload_verticalCompare = io_input_payload_verticalCompare;
  assign io_outputs_0_payload_mainDiff = io_input_payload_mainDiff;
  assign io_outputs_0_payload_counterDiff = io_input_payload_counterDiff;
  assign io_outputs_0_payload_horizontalDiff = io_input_payload_horizontalDiff;
  assign io_outputs_0_payload_verticalDiff = io_input_payload_verticalDiff;
  assign io_outputs_0_payload_isHorizontalMin = io_input_payload_isHorizontalMin;
  assign io_outputs_0_payload_minDiff = io_input_payload_minDiff;
  assign io_outputs_0_payload_currentPosition = io_input_payload_currentPosition;
  assign io_outputs_0_payload_nextPosition = io_input_payload_nextPosition;
  assign io_outputs_0_payload_horizontalDirectionValid = io_input_payload_horizontalDirectionValid;
  assign io_outputs_0_payload_verticalDirectionValid = io_input_payload_verticalDirectionValid;
  assign io_outputs_0_payload_mainDirectionValid = io_input_payload_mainDirectionValid;
  assign io_outputs_0_payload_counterDirectionValid = io_input_payload_counterDirectionValid;
  assign io_outputs_0_payload_inValidMinDiff = io_input_payload_inValidMinDiff;
  assign io_outputs_1_payload_frameStart = io_input_payload_frameStart;
  assign io_outputs_1_payload_rowEnd = io_input_payload_rowEnd;
  assign io_outputs_1_payload_pipeValid = io_input_payload_pipeValid;
  assign io_outputs_1_payload_firstRow = io_input_payload_firstRow;
  assign io_outputs_1_payload_lastRow = io_input_payload_lastRow;
  assign io_outputs_1_payload_finalResult = io_input_payload_finalResult;
  assign io_outputs_1_payload_mainCompare = io_input_payload_mainCompare;
  assign io_outputs_1_payload_counterCompare = io_input_payload_counterCompare;
  assign io_outputs_1_payload_horizontalCompare = io_input_payload_horizontalCompare;
  assign io_outputs_1_payload_verticalCompare = io_input_payload_verticalCompare;
  assign io_outputs_1_payload_mainDiff = io_input_payload_mainDiff;
  assign io_outputs_1_payload_counterDiff = io_input_payload_counterDiff;
  assign io_outputs_1_payload_horizontalDiff = io_input_payload_horizontalDiff;
  assign io_outputs_1_payload_verticalDiff = io_input_payload_verticalDiff;
  assign io_outputs_1_payload_isHorizontalMin = io_input_payload_isHorizontalMin;
  assign io_outputs_1_payload_minDiff = io_input_payload_minDiff;
  assign io_outputs_1_payload_currentPosition = io_input_payload_currentPosition;
  assign io_outputs_1_payload_nextPosition = io_input_payload_nextPosition;
  assign io_outputs_1_payload_horizontalDirectionValid = io_input_payload_horizontalDirectionValid;
  assign io_outputs_1_payload_verticalDirectionValid = io_input_payload_verticalDirectionValid;
  assign io_outputs_1_payload_mainDirectionValid = io_input_payload_mainDirectionValid;
  assign io_outputs_1_payload_counterDirectionValid = io_input_payload_counterDirectionValid;
  assign io_outputs_1_payload_inValidMinDiff = io_input_payload_inValidMinDiff;

endmodule

module StreamFork_2 (
  input               io_input_valid,
  output              io_input_ready,
  input               io_input_payload_frameStart,
  input               io_input_payload_rowEnd,
  input               io_input_payload_passMode,
  input               io_input_payload_passValid,
  input      [2:0]    io_input_payload_onceMode,
  input               io_input_payload_onceValid,
  input               io_input_payload_mainCompare,
  input               io_input_payload_counterCompare,
  input      [7:0]    io_input_payload_mainDiff,
  input      [7:0]    io_input_payload_counterDiff,
  input               io_input_payload_twiceCompValid,
  input      [2:0]    io_input_payload_twiceMode,
  input               io_input_payload_inpValidFlag,
  input               io_input_payload_oddValid,
  output              io_outputs_0_valid,
  input               io_outputs_0_ready,
  output              io_outputs_0_payload_frameStart,
  output              io_outputs_0_payload_rowEnd,
  output              io_outputs_0_payload_passMode,
  output              io_outputs_0_payload_passValid,
  output     [2:0]    io_outputs_0_payload_onceMode,
  output              io_outputs_0_payload_onceValid,
  output              io_outputs_0_payload_mainCompare,
  output              io_outputs_0_payload_counterCompare,
  output     [7:0]    io_outputs_0_payload_mainDiff,
  output     [7:0]    io_outputs_0_payload_counterDiff,
  output              io_outputs_0_payload_twiceCompValid,
  output     [2:0]    io_outputs_0_payload_twiceMode,
  output              io_outputs_0_payload_inpValidFlag,
  output              io_outputs_0_payload_oddValid,
  output              io_outputs_1_valid,
  input               io_outputs_1_ready,
  output              io_outputs_1_payload_frameStart,
  output              io_outputs_1_payload_rowEnd,
  output              io_outputs_1_payload_passMode,
  output              io_outputs_1_payload_passValid,
  output     [2:0]    io_outputs_1_payload_onceMode,
  output              io_outputs_1_payload_onceValid,
  output              io_outputs_1_payload_mainCompare,
  output              io_outputs_1_payload_counterCompare,
  output     [7:0]    io_outputs_1_payload_mainDiff,
  output     [7:0]    io_outputs_1_payload_counterDiff,
  output              io_outputs_1_payload_twiceCompValid,
  output     [2:0]    io_outputs_1_payload_twiceMode,
  output              io_outputs_1_payload_inpValidFlag,
  output              io_outputs_1_payload_oddValid
);


  assign io_input_ready = (io_outputs_0_ready && io_outputs_1_ready);
  assign io_outputs_0_valid = (io_input_valid && io_input_ready);
  assign io_outputs_1_valid = (io_input_valid && io_input_ready);
  assign io_outputs_0_payload_frameStart = io_input_payload_frameStart;
  assign io_outputs_0_payload_rowEnd = io_input_payload_rowEnd;
  assign io_outputs_0_payload_passMode = io_input_payload_passMode;
  assign io_outputs_0_payload_passValid = io_input_payload_passValid;
  assign io_outputs_0_payload_onceMode = io_input_payload_onceMode;
  assign io_outputs_0_payload_onceValid = io_input_payload_onceValid;
  assign io_outputs_0_payload_mainCompare = io_input_payload_mainCompare;
  assign io_outputs_0_payload_counterCompare = io_input_payload_counterCompare;
  assign io_outputs_0_payload_mainDiff = io_input_payload_mainDiff;
  assign io_outputs_0_payload_counterDiff = io_input_payload_counterDiff;
  assign io_outputs_0_payload_twiceCompValid = io_input_payload_twiceCompValid;
  assign io_outputs_0_payload_twiceMode = io_input_payload_twiceMode;
  assign io_outputs_0_payload_inpValidFlag = io_input_payload_inpValidFlag;
  assign io_outputs_0_payload_oddValid = io_input_payload_oddValid;
  assign io_outputs_1_payload_frameStart = io_input_payload_frameStart;
  assign io_outputs_1_payload_rowEnd = io_input_payload_rowEnd;
  assign io_outputs_1_payload_passMode = io_input_payload_passMode;
  assign io_outputs_1_payload_passValid = io_input_payload_passValid;
  assign io_outputs_1_payload_onceMode = io_input_payload_onceMode;
  assign io_outputs_1_payload_onceValid = io_input_payload_onceValid;
  assign io_outputs_1_payload_mainCompare = io_input_payload_mainCompare;
  assign io_outputs_1_payload_counterCompare = io_input_payload_counterCompare;
  assign io_outputs_1_payload_mainDiff = io_input_payload_mainDiff;
  assign io_outputs_1_payload_counterDiff = io_input_payload_counterDiff;
  assign io_outputs_1_payload_twiceCompValid = io_input_payload_twiceCompValid;
  assign io_outputs_1_payload_twiceMode = io_input_payload_twiceMode;
  assign io_outputs_1_payload_inpValidFlag = io_input_payload_inpValidFlag;
  assign io_outputs_1_payload_oddValid = io_input_payload_oddValid;

endmodule

module StreamFork_1 (
  input               io_input_valid,
  output              io_input_ready,
  input               io_input_payload_frameStart,
  input               io_input_payload_rowEnd,
  input               io_input_payload_passMode,
  input               io_input_payload_passValid,
  input      [2:0]    io_input_payload_onceMode,
  input               io_input_payload_onceValid,
  input               io_input_payload_mainCompare,
  input               io_input_payload_counterCompare,
  input      [7:0]    io_input_payload_mainDiff,
  input      [7:0]    io_input_payload_counterDiff,
  input               io_input_payload_twiceCompValid,
  input      [2:0]    io_input_payload_twiceMode,
  output              io_outputs_0_valid,
  input               io_outputs_0_ready,
  output              io_outputs_0_payload_frameStart,
  output              io_outputs_0_payload_rowEnd,
  output              io_outputs_0_payload_passMode,
  output              io_outputs_0_payload_passValid,
  output     [2:0]    io_outputs_0_payload_onceMode,
  output              io_outputs_0_payload_onceValid,
  output              io_outputs_0_payload_mainCompare,
  output              io_outputs_0_payload_counterCompare,
  output     [7:0]    io_outputs_0_payload_mainDiff,
  output     [7:0]    io_outputs_0_payload_counterDiff,
  output              io_outputs_0_payload_twiceCompValid,
  output     [2:0]    io_outputs_0_payload_twiceMode,
  output              io_outputs_1_valid,
  input               io_outputs_1_ready,
  output              io_outputs_1_payload_frameStart,
  output              io_outputs_1_payload_rowEnd,
  output              io_outputs_1_payload_passMode,
  output              io_outputs_1_payload_passValid,
  output     [2:0]    io_outputs_1_payload_onceMode,
  output              io_outputs_1_payload_onceValid,
  output              io_outputs_1_payload_mainCompare,
  output              io_outputs_1_payload_counterCompare,
  output     [7:0]    io_outputs_1_payload_mainDiff,
  output     [7:0]    io_outputs_1_payload_counterDiff,
  output              io_outputs_1_payload_twiceCompValid,
  output     [2:0]    io_outputs_1_payload_twiceMode
);


  assign io_input_ready = (io_outputs_0_ready && io_outputs_1_ready);
  assign io_outputs_0_valid = (io_input_valid && io_input_ready);
  assign io_outputs_1_valid = (io_input_valid && io_input_ready);
  assign io_outputs_0_payload_frameStart = io_input_payload_frameStart;
  assign io_outputs_0_payload_rowEnd = io_input_payload_rowEnd;
  assign io_outputs_0_payload_passMode = io_input_payload_passMode;
  assign io_outputs_0_payload_passValid = io_input_payload_passValid;
  assign io_outputs_0_payload_onceMode = io_input_payload_onceMode;
  assign io_outputs_0_payload_onceValid = io_input_payload_onceValid;
  assign io_outputs_0_payload_mainCompare = io_input_payload_mainCompare;
  assign io_outputs_0_payload_counterCompare = io_input_payload_counterCompare;
  assign io_outputs_0_payload_mainDiff = io_input_payload_mainDiff;
  assign io_outputs_0_payload_counterDiff = io_input_payload_counterDiff;
  assign io_outputs_0_payload_twiceCompValid = io_input_payload_twiceCompValid;
  assign io_outputs_0_payload_twiceMode = io_input_payload_twiceMode;
  assign io_outputs_1_payload_frameStart = io_input_payload_frameStart;
  assign io_outputs_1_payload_rowEnd = io_input_payload_rowEnd;
  assign io_outputs_1_payload_passMode = io_input_payload_passMode;
  assign io_outputs_1_payload_passValid = io_input_payload_passValid;
  assign io_outputs_1_payload_onceMode = io_input_payload_onceMode;
  assign io_outputs_1_payload_onceValid = io_input_payload_onceValid;
  assign io_outputs_1_payload_mainCompare = io_input_payload_mainCompare;
  assign io_outputs_1_payload_counterCompare = io_input_payload_counterCompare;
  assign io_outputs_1_payload_mainDiff = io_input_payload_mainDiff;
  assign io_outputs_1_payload_counterDiff = io_input_payload_counterDiff;
  assign io_outputs_1_payload_twiceCompValid = io_input_payload_twiceCompValid;
  assign io_outputs_1_payload_twiceMode = io_input_payload_twiceMode;

endmodule

module StreamFork (
  input               io_input_valid,
  output              io_input_ready,
  input      [31:0]   io_input_payload_pixel,
  input               io_input_payload_frameStart,
  input               io_input_payload_rowEnd,
  output              io_outputs_0_valid,
  input               io_outputs_0_ready,
  output     [31:0]   io_outputs_0_payload_pixel,
  output              io_outputs_0_payload_frameStart,
  output              io_outputs_0_payload_rowEnd,
  output              io_outputs_1_valid,
  input               io_outputs_1_ready,
  output     [31:0]   io_outputs_1_payload_pixel,
  output              io_outputs_1_payload_frameStart,
  output              io_outputs_1_payload_rowEnd,
  output              io_outputs_2_valid,
  input               io_outputs_2_ready,
  output     [31:0]   io_outputs_2_payload_pixel,
  output              io_outputs_2_payload_frameStart,
  output              io_outputs_2_payload_rowEnd
);


  assign io_input_ready = ((io_outputs_0_ready && io_outputs_1_ready) && io_outputs_2_ready);
  assign io_outputs_0_valid = (io_input_valid && io_input_ready);
  assign io_outputs_1_valid = (io_input_valid && io_input_ready);
  assign io_outputs_2_valid = (io_input_valid && io_input_ready);
  assign io_outputs_0_payload_pixel = io_input_payload_pixel;
  assign io_outputs_0_payload_frameStart = io_input_payload_frameStart;
  assign io_outputs_0_payload_rowEnd = io_input_payload_rowEnd;
  assign io_outputs_1_payload_pixel = io_input_payload_pixel;
  assign io_outputs_1_payload_frameStart = io_input_payload_frameStart;
  assign io_outputs_1_payload_rowEnd = io_input_payload_rowEnd;
  assign io_outputs_2_payload_pixel = io_input_payload_pixel;
  assign io_outputs_2_payload_frameStart = io_input_payload_frameStart;
  assign io_outputs_2_payload_rowEnd = io_input_payload_rowEnd;

endmodule

module StreamTransactionCounter (
  input               io_ctrlFire,
  input               io_targetFire,
  input      [9:0]    io_count,
  output              io_working,
  output              io_last,
  output              io_done,
  output     [9:0]    io_value,
  input               clk,
  input               resetn
);

  wire       [9:0]    CICC1851_counter_valueNext;
  wire       [0:0]    CICC1851_counter_valueNext_1;
  reg        [9:0]    countReg;
  reg                 counter_willIncrement;
  reg                 counter_willClear;
  reg        [9:0]    counter_valueNext;
  reg        [9:0]    counter_value;
  wire                counter_willOverflowIfInc;
  wire                counter_willOverflow;
  wire       [9:0]    expected;
  wire                lastOne;
  reg                 running;
  wire                done;
  wire                doneWithFire;
  wire                when_Stream_l1776;

  assign CICC1851_counter_valueNext_1 = counter_willIncrement;
  assign CICC1851_counter_valueNext = {9'd0, CICC1851_counter_valueNext_1};
  always @(*) begin
    counter_willIncrement = 1'b0;
    if(!done) begin
      if(io_targetFire) begin
        counter_willIncrement = 1'b1;
      end
    end
  end

  always @(*) begin
    counter_willClear = 1'b0;
    if(done) begin
      counter_willClear = 1'b1;
    end
  end

  assign counter_willOverflowIfInc = (counter_value == 10'h3ff);
  assign counter_willOverflow = (counter_willOverflowIfInc && counter_willIncrement);
  always @(*) begin
    counter_valueNext = (counter_value + CICC1851_counter_valueNext);
    if(counter_willClear) begin
      counter_valueNext = 10'h0;
    end
  end

  assign expected = countReg;
  assign lastOne = (counter_value == expected);
  assign done = (lastOne && io_targetFire);
  assign doneWithFire = 1'b1;
  assign when_Stream_l1776 = (done && io_ctrlFire);
  assign io_working = running;
  assign io_last = lastOne;
  assign io_done = (lastOne && io_targetFire);
  assign io_value = counter_value;
  always @(posedge clk) begin
    if(io_ctrlFire) begin
      countReg <= io_count;
    end
  end

  always @(posedge clk or negedge resetn) begin
    if(!resetn) begin
      counter_value <= 10'h0;
      running <= 1'b0;
    end else begin
      counter_value <= counter_valueNext;
      if(when_Stream_l1776) begin
        running <= doneWithFire;
      end else begin
        if(io_ctrlFire) begin
          running <= 1'b1;
        end else begin
          if(done) begin
            running <= 1'b0;
          end
        end
      end
    end
  end


endmodule
